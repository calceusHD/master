library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity grng_pwclt12 is port(
  iClk : in std_logic;
  iCE : in std_logic := '1';
  iLoadEn : in std_logic := '0';
  iLoadData : in std_logic := '0';
  oRes : out std_logic_vector(26-1 downto 0)
); end entity;

architecture RTL of grng_pwclt12 is
    signal iURNG : std_logic_vector(300-1 downto 0);
    --Bernoulli
    -- bernoulli_fp, fb=52, frac_width=51, exp_width=7
    --   exp_src_width=119
    signal bernoulli_fp_out : boolean;
    signal bernoulli_fp_thresh : unsigned(58-1 downto 0);
    signal bernoulli_fp_urng : std_logic_vector(170-1 downto 0);
    signal bernoulli_fp_cx_exp_urng : std_logic_vector(119-1 downto 0);
    signal bernoulli_fp_c0_frac_thresh, bernoulli_fp_c0_frac_rand : unsigned(51-1 downto 0);
    signal bernoulli_fp_cx_exp_rand, bernoulli_fp_c0_exp_thresh: unsigned(7-1 downto 0);
    signal bernoulli_fp_c1_exp_greater, bernoulli_fp_c1_exp_equal, bernoulli_fp_c1_frac_greater : boolean;
    signal lmz_branch_1, lmz_branch_1_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_1, lmz_branch_hit_1_sig : boolean;
    signal lmz_branch_2, lmz_branch_2_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_2, lmz_branch_hit_2_sig : boolean;
    signal lmz_branch_3, lmz_branch_3_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_3, lmz_branch_hit_3_sig : boolean;
    signal lmz_branch_4, lmz_branch_4_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_4, lmz_branch_hit_4_sig : boolean;
    signal lmz_branch_5, lmz_branch_5_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_5, lmz_branch_hit_5_sig : boolean;
    signal lmz_branch_6, lmz_branch_6_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_6, lmz_branch_hit_6_sig : boolean;
    signal lmz_branch_7, lmz_branch_7_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_7, lmz_branch_hit_7_sig : boolean;
    signal lmz_branch_8, lmz_branch_8_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_8, lmz_branch_hit_8_sig : boolean;
    signal lmz_branch_9, lmz_branch_9_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_9, lmz_branch_hit_9_sig : boolean;
    signal lmz_branch_10, lmz_branch_10_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_10, lmz_branch_hit_10_sig : boolean;
    signal lmz_branch_11, lmz_branch_11_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_11, lmz_branch_hit_11_sig : boolean;
    signal lmz_branch_12, lmz_branch_12_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_12, lmz_branch_hit_12_sig : boolean;
    signal lmz_branch_13, lmz_branch_13_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_13, lmz_branch_hit_13_sig : boolean;
    signal lmz_branch_14, lmz_branch_14_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_14, lmz_branch_hit_14_sig : boolean;
    signal lmz_branch_15, lmz_branch_15_sig : unsigned(7-1 downto 0);
    signal lmz_branch_hit_15, lmz_branch_hit_15_sig : boolean;
    signal bernoulli_fp_c0_exp_rand : unsigned(7-1 downto 0);
    signal bernoulli_fp_c0_exp_rand_d1 : unsigned(7-1 downto 0);
    signal bernoulli_fp_c0_exp_rand_d2 : unsigned(7-1 downto 0);
    --Alias table
    signal alias_table_urng : std_logic_vector(179-1 downto 0);
    signal alias_table_out, c0_alias_index : unsigned(9-1 downto 0);
    attribute rom_style : string;
    type alias_rom_t is array(0 to 2*512-1) of unsigned(34-1 downto 0);
    signal alias_rom : alias_rom_t := (
        "0000101110111110100011100000111100", -- i=0, alt=60, thresh=0.983859, actual=0.012471, err=0
        "0001000000000010111001111000001001", -- i=1, alt=9, thresh=0.811589, actual=0.0249298, err=0
        "0001011010111101001111101000101011", -- i=2, alt=43, thresh=0.817009, actual=0.0248933, err=-3.46945e-018
        "0110111111000010110111110000010101", -- i=3, alt=21, thresh=0.810736, actual=0.0248326, err=0
        "0000101000001100110010010001000100", -- i=4, alt=68, thresh=0.799622, actual=0.0247478, err=0
        "0100011110001110001110110000111011", -- i=5, alt=59, thresh=0.801928, actual=0.0246392, err=0
        "0110100001010011100011101000011110", -- i=6, alt=30, thresh=0.814068, actual=0.0245071, err=0
        "0111011000011011111001011000010110", -- i=7, alt=22, thresh=0.909361, actual=0.024352, err=-3.46945e-018
        "0001100000111000001101001000011001", -- i=8, alt=25, thresh=0.979439, actual=0.0241741, err=3.46945e-018
        "0001001111110111000000111000011001", -- i=9, alt=25, thresh=0.995288, actual=0.0239742, err=0
        "0110111101110010111000011000110101", -- i=10, alt=53, thresh=0.98305, actual=0.0237526, err=0
        "0011011000111111100010101000100010", -- i=11, alt=34, thresh=0.99903, actual=0.0235102, err=0
        "0111010110110110001110111000010000", -- i=12, alt=16, thresh=0.925006, actual=0.0232474, err=0
        "0011101111010110011101010000011010", -- i=13, alt=26, thresh=0.816642, actual=0.0229652, err=3.46945e-018
        "0111110101001100111010110000110000", -- i=14, alt=48, thresh=0.827525, actual=0.0226642, err=0
        "0100110010011111010100011000111100", -- i=15, alt=60, thresh=0.999979, actual=0.0223454, err=0
        "0010111011100000110100011000110101", -- i=16, alt=53, thresh=0.998163, actual=0.0220095, err=0
        "0101001010111101011000111001000011", -- i=17, alt=67, thresh=0.97289, actual=0.0216574, err=0
        "0111111001101111000011111000111101", -- i=18, alt=61, thresh=0.925519, actual=0.0212902, err=0
        "0000110111001011111001001000001000", -- i=19, alt=8, thresh=0.822349, actual=0.0209088, err=0
        "0110000001100011110110101000010101", -- i=20, alt=21, thresh=0.877578, actual=0.0205141, err=0
        "0101000010010011111100001000011110", -- i=21, alt=30, thresh=0.984397, actual=0.0201073, err=0
        "0011111110000111110100101000100011", -- i=22, alt=35, thresh=0.995708, actual=0.0196892, err=0
        "0101110011010001001100101001000111", -- i=23, alt=71, thresh=0.889482, actual=0.019261, err=-3.46945e-018
        "0111111000010000101011011000001000", -- i=24, alt=8, thresh=0.779261, actual=0.0188238, err=0
        "0100011001100011011010101000111101", -- i=25, alt=61, thresh=0.999696, actual=0.0183785, err=-3.46945e-018
        "0010100100100100100010000000100010", -- i=26, alt=34, thresh=0.997746, actual=0.0179261, err=0
        "0011101001111111011100100000011001", -- i=27, alt=25, thresh=0.961385, actual=0.0174679, err=0
        "0100100111001001001000001001000101", -- i=28, alt=69, thresh=0.812733, actual=0.0170047, err=0
        "0110110100001011101000100001001000", -- i=29, alt=72, thresh=0.985168, actual=0.0165377, err=0
        "0110110101100101100111001000001111", -- i=30, alt=15, thresh=0.998988, actual=0.0160678, err=0
        "0011001111000010001101001001000101", -- i=31, alt=69, thresh=0.99635, actual=0.0155959, err=-1.73472e-018
        "0100101010001100000010100000000000", -- i=32, alt=0, thresh=0.822242, actual=0.0151232, err=1.73472e-018
        "0101010110101001110110001000001001", -- i=33, alt=9, thresh=0.907593, actual=0.0146504, err=1.73472e-018
        "0101010110101001110110001000100010", -- i=34, alt=34, thresh=NaN, actual=0.0141786, err=-7.45931e-017
        "0100000101101110100101101000111100", -- i=35, alt=60, thresh=0.999133, actual=0.0137085, err=1.73472e-018
        "0110010001011111110001101000001010", -- i=36, alt=10, thresh=0.817939, actual=0.0132411, err=-1.73472e-018
        "0011110101110011111111101000111011", -- i=37, alt=59, thresh=0.83241, actual=0.0127772, err=0
        "0000001010000001111101011000001011", -- i=38, alt=11, thresh=0.985942, actual=0.0123174, err=0
        "0011111011010000101000010001000011", -- i=39, alt=67, thresh=0.998024, actual=0.0118626, err=-1.73472e-018
        "0000011011101111100011100000110100", -- i=40, alt=52, thresh=0.874731, actual=0.0114135, err=0
        "0000111101011011010100110000101111", -- i=41, alt=47, thresh=0.787299, actual=0.0109706, err=0
        "0110101100101000111011101000100111", -- i=42, alt=39, thresh=0.981144, actual=0.0105346, err=-3.46945e-018
        "0100000000000000000111101000111101", -- i=43, alt=61, thresh=0.994615, actual=0.010106, err=-1.73472e-018
        "0010100001000000001011100000011110", -- i=44, alt=30, thresh=0.971581, actual=0.00968546, err=0
        "0110011010110110010100010000100010", -- i=45, alt=34, thresh=0.812673, actual=0.00927331, err=0
        "0010111111101011001110111001000100", -- i=46, alt=68, thresh=0.857883, actual=0.00887002, err=-1.73472e-018
        "0100001001001000110110100000100111", -- i=47, alt=39, thresh=0.992082, actual=0.00847599, err=0
        "0111100101110101110110110000100011", -- i=48, alt=35, thresh=0.974662, actual=0.00809155, err=1.73472e-018
        "0111010101111101010010011000001011", -- i=49, alt=11, thresh=0.967011, actual=0.00771701, err=0
        "0000101100111000011110010000100110", -- i=50, alt=38, thresh=0.807314, actual=0.00735261, err=8.67362e-019
        "0101101101101011010000111000101010", -- i=51, alt=42, thresh=0.827372, actual=0.00699858, err=0
        "0111011100010010110010010000110110", -- i=52, alt=54, thresh=0.987416, actual=0.00665508, err=-8.67362e-019
        "0100001010000100101000101000100010", -- i=53, alt=34, thresh=0.999989, actual=0.00632227, err=0
        "0110010000010001111010101000001111", -- i=54, alt=15, thresh=0.999886, actual=0.00600023, err=-8.67362e-019
        "0101001111001010001000111000110110", -- i=55, alt=54, thresh=0.932737, actual=0.00568903, err=0
        "0101101111010100010110101000010000", -- i=56, alt=16, thresh=0.811748, actual=0.00538871, err=0
        "0010111111110010111011111000111100", -- i=57, alt=60, thresh=0.815139, actual=0.00509925, err=0
        "0110000100010010110111100000100010", -- i=58, alt=34, thresh=0.946377, actual=0.00482063, err=8.67362e-019
        "0011101010000101011110001001000101", -- i=59, alt=69, thresh=0.96625, actual=0.00455279, err=8.67362e-019
        "0101010100111101100110011000100010", -- i=60, alt=34, thresh=0.999996, actual=0.00429562, err=0
        "0010001111100001011111111001000011", -- i=61, alt=67, thresh=0.999904, actual=0.00404902, err=0
        "0110110011010101001110011000110101", -- i=62, alt=53, thresh=0.966358, actual=0.00381285, err=0
        "0010111110101001111000111000100110", -- i=63, alt=38, thresh=0.871084, actual=0.00358695, err=-4.33681e-019
        "0110101101010110100101111000110101", -- i=64, alt=53, thresh=0.813439, actual=0.00337114, err=0
        "0101100011101111111001010000000000", -- i=65, alt=0, thresh=0.775877, actual=0.00316522, err=0
        "0000001110101000010100000000101111", -- i=66, alt=47, thresh=0.864304, actual=0.00296897, err=0
        "0001101100100110011111101000111100", -- i=67, alt=60, thresh=0.999965, actual=0.00278217, err=0
        "0101110010100011100110111000010000", -- i=68, alt=16, thresh=0.991049, actual=0.00260458, err=-4.33681e-019
        "0001101101110001010011101000110110", -- i=69, alt=54, thresh=0.999746, actual=0.00243594, err=-4.33681e-019
        "0101001100111100010110110000100010", -- i=70, alt=34, thresh=0.983018, actual=0.00227599, err=0
        "0010111100111101111000010001000101", -- i=71, alt=69, thresh=0.977213, actual=0.00212447, err=0
        "0111010111010010111011001001000011", -- i=72, alt=67, thresh=0.999494, actual=0.0019811, err=0
        "0101000111001111100101001000100111", -- i=73, alt=39, thresh=0.94495, actual=0.00184561, err=2.1684e-019
        "0010111100000010010001101000010001", -- i=74, alt=17, thresh=0.87946, actual=0.0017177, err=2.1684e-019
        "0000100001111011100000110001000110", -- i=75, alt=70, thresh=0.817709, actual=0.00159709, err=2.1684e-019
        "0110101101101000011100101000101010", -- i=76, alt=42, thresh=0.759552, actual=0.0014835, err=0
        "0101010101110010000110111000110100", -- i=77, alt=52, thresh=0.704841, actual=0.00137664, err=0
        "0001100111000111010100111000011001", -- i=78, alt=25, thresh=0.653433, actual=0.00127624, err=0
        "0110001000010100101011110001000011", -- i=79, alt=67, thresh=0.605182, actual=0.001182, err=2.1684e-019
        "0100010000011010110100110000001111", -- i=80, alt=15, thresh=0.559947, actual=0.00109365, err=2.1684e-019
        "0101101110110100000110100000011101", -- i=81, alt=29, thresh=0.517587, actual=0.00101091, err=0
        "0010000111111111010011001000111010", -- i=82, alt=58, thresh=0.477964, actual=0.000933524, err=0
        "0101011000101010011111000000000111", -- i=83, alt=7, thresh=0.440944, actual=0.000861218, err=1.0842e-019
        "0001001000110110010110110000100001", -- i=84, alt=33, thresh=0.406393, actual=0.000793737, err=0
        "0010101110101010100101000000010100", -- i=85, alt=20, thresh=0.374184, actual=0.000730828, err=1.0842e-019
        "0000100110001110011001111001000010", -- i=86, alt=66, thresh=0.344191, actual=0.000672249, err=0
        "0100011110001111001110110000101110", -- i=87, alt=46, thresh=0.316293, actual=0.00061776, err=0
        "0001000011000010000111110000100101", -- i=88, alt=37, thresh=0.290373, actual=0.000567134, err=1.0842e-019
        "0011101100011101101111011000000110", -- i=89, alt=6, thresh=0.266316, actual=0.000520148, err=0
        "0101000100001011100111101000110011", -- i=90, alt=51, thresh=0.244014, actual=0.000476589, err=0
        "0101111010000010100111010000001110", -- i=91, alt=14, thresh=0.223361, actual=0.000436251, err=5.42101e-020
        "0001001111001010011100110000111001", -- i=92, alt=57, thresh=0.204256, actual=0.000398937, err=5.42101e-020
        "0001110000010011010111011000000101", -- i=93, alt=5, thresh=0.186603, actual=0.000364459, err=5.42101e-020
        "0101001011100001001011010000101001", -- i=94, alt=41, thresh=0.170309, actual=0.000332635, err=0
        "0100110100001001100001111001000001", -- i=95, alt=65, thresh=0.155286, actual=0.000303293, err=0
        "0111011001100000011101001000011000", -- i=96, alt=24, thresh=0.14145, actual=0.00027627, err=0
        "0100111111000000011111010000000100", -- i=97, alt=4, thresh=0.128721, actual=0.000251408, err=5.42101e-020
        "0100000001000000000001011000010011", -- i=98, alt=19, thresh=0.117023, actual=0.00022856, err=0
        "0110011100011111010000010000011100", -- i=99, alt=28, thresh=0.106284, actual=0.000207586, err=0
        "0001100001000111000101000000000011", -- i=100, alt=3, thresh=0.0964365, actual=0.000188353, err=2.71051e-020
        "0110010110000000100110011001000000", -- i=101, alt=64, thresh=0.0874158, actual=0.000170734, err=0
        "0100000011000101100100111000100000", -- i=102, alt=32, thresh=0.0791616, actual=0.000154612, err=0
        "0000011100111010111101100000000010", -- i=103, alt=2, thresh=0.0716167, actual=0.000139876, err=2.71051e-020
        "0110001100001010100010101000101101", -- i=104, alt=45, thresh=0.0647276, actual=0.000126421, err=2.71051e-020
        "0111010000011010010001010000001101", -- i=105, alt=13, thresh=0.0584441, actual=0.000114149, err=1.35525e-020
        "0110110111011100000100110000111000", -- i=106, alt=56, thresh=0.052719, actual=0.000102967, err=0
        "0010010001011100010011101000000001", -- i=107, alt=1, thresh=0.0475083, actual=9.27897e-005, err=1.35525e-020
        "0010111111110011111010110000110010", -- i=108, alt=50, thresh=0.0427708, actual=8.35367e-005, err=0
        "0111110111101101111111011000100100", -- i=109, alt=36, thresh=0.0384681, actual=7.5133e-005, err=1.35525e-020
        "0111010110110001010001010000111111", -- i=110, alt=63, thresh=0.0345645, actual=6.75087e-005, err=1.35525e-020
        "0010111000111100101100101000101000", -- i=111, alt=40, thresh=0.0310266, actual=6.05989e-005, err=6.77626e-021
        "0111110010000000001111010000010111", -- i=112, alt=23, thresh=0.0278237, actual=5.43432e-005, err=0
        "0100001001001000100001010000010010", -- i=113, alt=18, thresh=0.024927, actual=4.86856e-005, err=0
        "0000011011111101011000000000001100", -- i=114, alt=12, thresh=0.0223101, actual=4.35745e-005, err=6.77626e-021
        "0000000011111011011110011000110111", -- i=115, alt=55, thresh=0.0199485, actual=3.89618e-005, err=0
        "0101101110101000001011001000011011", -- i=116, alt=27, thresh=0.0178194, actual=3.48034e-005, err=6.77626e-021
        "0111011011010000000000101000110001", -- i=117, alt=49, thresh=0.015902, actual=3.10585e-005, err=6.77626e-021
        "0100010100001111100000000000111110", -- i=118, alt=62, thresh=0.014177, actual=2.76895e-005, err=0
        "0010010100110111101001011000101100", -- i=119, alt=44, thresh=0.0126268, actual=2.46618e-005, err=3.38813e-021
        "0110111111011011101101011000011111", -- i=120, alt=31, thresh=0.0112352, actual=2.19437e-005, err=0
        "0011101000000100000111110000100011", -- i=121, alt=35, thresh=0.00998711, actual=1.95061e-005, err=3.38813e-021
        "0001101100001010110011111000001011", -- i=122, alt=11, thresh=0.00886903, actual=1.73223e-005, err=3.38813e-021
        "0110110111000010011100001000110110", -- i=123, alt=54, thresh=0.00786843, actual=1.5368e-005, err=0
        "0100100010011001110100010000111101", -- i=124, alt=61, thresh=0.0069739, actual=1.36209e-005, err=1.69407e-021
        "0001011110010101110101010000100111", -- i=125, alt=39, thresh=0.00617503, actual=1.20606e-005, err=1.69407e-021
        "0010010001011001101111110000010110", -- i=126, alt=22, thresh=0.00546233, actual=1.06686e-005, err=1.69407e-021
        "0001110011110110001000101000010001", -- i=127, alt=17, thresh=0.00482717, actual=9.42806e-006, err=1.69407e-021
        "0110011010100110100011110000110000", -- i=128, alt=48, thresh=0.0042617, actual=8.32362e-006, err=1.69407e-021
        "0101001000101011110110001000001010", -- i=129, alt=10, thresh=0.00375879, actual=7.34139e-006, err=8.47033e-022
        "0001000100111111101110001000101011", -- i=130, alt=43, thresh=0.00331199, actual=6.46873e-006, err=8.47033e-022
        "0000100011011011001101101000011010", -- i=131, alt=26, thresh=0.00291545, actual=5.69424e-006, err=8.47033e-022
        "0001111101011101000000001000111100", -- i=132, alt=60, thresh=0.00256389, actual=5.00759e-006, err=8.47033e-022
        "0010110101000011001100100000011110", -- i=133, alt=30, thresh=0.00225251, actual=4.39943e-006, err=0
        "0110001100010001100001001000110101", -- i=134, alt=53, thresh=0.00197702, actual=3.86136e-006, err=8.47033e-022
        "0100011011111000100101010000100010", -- i=135, alt=34, thresh=0.00173352, actual=3.38579e-006, err=4.23516e-022
        "0110001100111011000100111000010000", -- i=136, alt=16, thresh=0.00151853, actual=2.96589e-006, err=4.23516e-022
        "0001110110111000110001010000001001", -- i=137, alt=9, thresh=0.00132891, actual=2.59552e-006, err=0
        "0010110000100100101010000000010101", -- i=138, alt=21, thresh=0.00116183, actual=2.26919e-006, err=4.23516e-022
        "0001010101100100000111111000100110", -- i=139, alt=38, thresh=0.00101476, actual=1.98195e-006, err=4.23516e-022
        "0101001000010101010000110000111011", -- i=140, alt=59, thresh=0.000885442, actual=1.72938e-006, err=0
        "0111000010101110000110111000101111", -- i=141, alt=47, thresh=0.00077185, actual=1.50752e-006, err=2.11758e-022
        "0100101111000001101100110000001000", -- i=142, alt=8, thresh=0.000672174, actual=1.31284e-006, err=0
        "0000101101010000011000110000000000", -- i=143, alt=0, thresh=0.000584798, actual=1.14218e-006, err=2.11758e-022
        "0100101001111010111001101000101010", -- i=144, alt=42, thresh=0.000508283, actual=9.9274e-007, err=2.11758e-022
        "0011001101001000111001110000110100", -- i=145, alt=52, thresh=0.000441348, actual=8.62007e-007, err=0
        "0111111011110000000111000000011001", -- i=146, alt=25, thresh=0.000382853, actual=7.47759e-007, err=0
        "0101101000110010100100011000001111", -- i=147, alt=15, thresh=0.000331786, actual=6.4802e-007, err=1.05879e-022
        "0111111001000100101100010000011101", -- i=148, alt=29, thresh=0.00028725, actual=5.61036e-007, err=1.05879e-022
        "0001010100101010000110000000111010", -- i=149, alt=58, thresh=0.00024845, actual=4.85253e-007, err=0
        "0111000101011001010110100000000111", -- i=150, alt=7, thresh=0.00021468, actual=4.19297e-007, err=5.29396e-023
        "0111001011000100101011100000100001", -- i=151, alt=33, thresh=0.000185319, actual=3.61952e-007, err=5.29396e-023
        "0101111111110011000000011000010100", -- i=152, alt=20, thresh=0.000159818, actual=3.12144e-007, err=5.29396e-023
        "0000101110111001001010101000101110", -- i=153, alt=46, thresh=0.000137691, actual=2.68928e-007, err=5.29396e-023
        "0110100110100101010010110000100101", -- i=154, alt=37, thresh=0.000118512, actual=2.31468e-007, err=0
        "0100001101111001011011110000000110", -- i=155, alt=6, thresh=0.000101904, actual=1.99032e-007, err=2.64698e-023
        "0010011100111000110110011000110011", -- i=156, alt=51, thresh=8.75387e-005, actual=1.70974e-007, err=2.64698e-023
        "0100100010000100000011100000001110", -- i=157, alt=14, thresh=7.51247e-005, actual=1.46728e-007, err=2.64698e-023
        "0010011111100110110100001000111001", -- i=158, alt=57, thresh=6.44082e-005, actual=1.25797e-007, err=2.64698e-023
        "0111101111001110100101100000000101", -- i=159, alt=5, thresh=5.51664e-005, actual=1.07747e-007, err=1.32349e-023
        "0010001111000000001101101000101001", -- i=160, alt=41, thresh=4.72046e-005, actual=9.21965e-008, err=1.32349e-023
        "0001010110100011110110110000011000", -- i=161, alt=24, thresh=4.03524e-005, actual=7.88133e-008, err=1.32349e-023
        "0111110110001110111101101000000100", -- i=162, alt=4, thresh=3.44612e-005, actual=6.7307e-008, err=0
        "0111110000000111100111100000010011", -- i=163, alt=19, thresh=2.94013e-005, actual=5.74244e-008, err=0
        "0110100001111100000111000000011100", -- i=164, alt=28, thresh=2.50598e-005, actual=4.8945e-008, err=6.61744e-024
        "0001111010010100100000001000000011", -- i=165, alt=3, thresh=2.13386e-005, actual=4.1677e-008, err=6.61744e-024
        "0001110111001111010111101000100000", -- i=166, alt=32, thresh=1.81522e-005, actual=3.54535e-008, err=0
        "0100001111000000100111110000000010", -- i=167, alt=2, thresh=1.54265e-005, actual=3.01299e-008, err=6.61744e-024
        "0011010011100011100111010000101101", -- i=168, alt=45, thresh=1.30973e-005, actual=2.55807e-008, err=3.30872e-024
        "0000001011000011101001001000001101", -- i=169, alt=13, thresh=1.11089e-005, actual=2.16971e-008, err=0
        "0110111011011000001000001000111000", -- i=170, alt=56, thresh=9.41321e-006, actual=1.83852e-008, err=0
        "0000100110001111001010011000000001", -- i=171, alt=1, thresh=7.96854e-006, actual=1.55636e-008, err=0
        "0011010011001101011111110000110010", -- i=172, alt=50, thresh=6.739e-006, actual=1.31621e-008, err=0
        "0111111101111001101100000000100100", -- i=173, alt=36, thresh=5.69362e-006, actual=1.11203e-008, err=1.65436e-024
        "0000010111111010100010110000101000", -- i=174, alt=40, thresh=4.80569e-006, actual=9.38612e-009, err=1.65436e-024
        "0000101000010011000001110000010111", -- i=175, alt=23, thresh=4.05228e-006, actual=7.91462e-009, err=1.65436e-024
        "0110011110111000111010110000010010", -- i=176, alt=18, thresh=3.41365e-006, actual=6.66729e-009, err=8.27181e-025
        "0100100110010101111000001000001100", -- i=177, alt=12, thresh=2.87286e-006, actual=5.61105e-009, err=0
        "0110100001111001101111001000110111", -- i=178, alt=55, thresh=2.41537e-006, actual=4.71753e-009, err=8.27181e-025
        "0010010001111000000000111000011011", -- i=179, alt=27, thresh=2.02876e-006, actual=3.96242e-009, err=0
        "0101110010110101000111111000110001", -- i=180, alt=49, thresh=1.70236e-006, actual=3.32493e-009, err=0
        "0011000100011111111000010000101100", -- i=181, alt=44, thresh=1.42708e-006, actual=2.78727e-009, err=4.1359e-025
        "0110100111010000110001011000011111", -- i=182, alt=31, thresh=1.19515e-006, actual=2.33428e-009, err=4.1359e-025
        "0011110100100000101111010000100011", -- i=183, alt=35, thresh=9.99932e-007, actual=1.95299e-009, err=0
        "0111111011101100011000001000001011", -- i=184, alt=11, thresh=8.35785e-007, actual=1.63239e-009, err=0
        "0011010100010011111111110000110110", -- i=185, alt=54, thresh=6.97902e-007, actual=1.36309e-009, err=0
        "0010101110101100101000010000100111", -- i=186, alt=39, thresh=5.82197e-007, actual=1.1371e-009, err=2.06795e-025
        "0001101011100001000000000000010110", -- i=187, alt=22, thresh=4.852e-007, actual=9.47656e-010, err=2.06795e-025
        "0001110001000101111001100000010001", -- i=188, alt=17, thresh=4.03968e-007, actual=7.89e-010, err=0
        "0110111000010010001110011000110000", -- i=189, alt=48, thresh=3.36008e-007, actual=6.56265e-010, err=1.03398e-025
        "0001001001110111011111000000001010", -- i=190, alt=10, thresh=2.79207e-007, actual=5.45327e-010, err=0
        "0001001011101001001111011000101011", -- i=191, alt=43, thresh=2.31782e-007, actual=4.527e-010, err=0
        "0111101110101011011011100000011010", -- i=192, alt=26, thresh=1.92225e-007, actual=3.75439e-010, err=0
        "0010101111000000101000110000011110", -- i=193, alt=30, thresh=1.59263e-007, actual=3.1106e-010, err=0
        "0111101010101010101011010000110101", -- i=194, alt=53, thresh=1.31824e-007, actual=2.57469e-010, err=0
        "0101111111000010011100011000100010", -- i=195, alt=34, thresh=1.09006e-007, actual=2.12902e-010, err=0
        "0010110000111100111010001000010000", -- i=196, alt=16, thresh=9.00495e-008, actual=1.75878e-010, err=0
        "0101101011010111101000111000001001", -- i=197, alt=9, thresh=7.4317e-008, actual=1.4515e-010, err=0
        "0101011111011110001100010000010101", -- i=198, alt=21, thresh=6.12732e-008, actual=1.19674e-010, err=0
        "0110011101110010011111101000100110", -- i=199, alt=38, thresh=5.04695e-008, actual=9.85733e-011, err=1.29247e-026
        "0101001001111001111011101000101111", -- i=200, alt=47, thresh=4.15301e-008, actual=8.11135e-011, err=1.29247e-026
        "0000101001110011010101000000001000", -- i=201, alt=8, thresh=3.41407e-008, actual=6.6681e-011, err=0
        "0100010110001001110010011000000000", -- i=202, alt=0, thresh=2.80387e-008, actual=5.4763e-011, err=6.46235e-027
        "0000100100001111011010111000101010", -- i=203, alt=42, thresh=2.30048e-008, actual=4.49312e-011, err=6.46235e-027
        "0010111001011101010101111000110100", -- i=204, alt=52, thresh=1.88562e-008, actual=3.68285e-011, err=6.46235e-027
        "0110011110001001000101110000011001", -- i=205, alt=25, thresh=1.54407e-008, actual=3.01576e-011, err=6.46235e-027
        "0111000001100111000101011000001111", -- i=206, alt=15, thresh=1.26315e-008, actual=2.46708e-011, err=3.23117e-027
        "0011011110000101110000101000011101", -- i=207, alt=29, thresh=1.03233e-008, actual=2.01626e-011, err=3.23117e-027
        "0100001101000100011111010000000111", -- i=208, alt=7, thresh=8.4286e-009, actual=1.64621e-011, err=0
        "0010111001000000001011011000100001", -- i=209, alt=33, thresh=6.87495e-009, actual=1.34276e-011, err=0
        "0100110101000111010001000000010100", -- i=210, alt=20, thresh=5.60221e-009, actual=1.09418e-011, err=0
        "0000111001111010001101001000101110", -- i=211, alt=46, thresh=4.56063e-009, actual=8.90749e-012, err=1.61559e-027
        "0010101100000001011111011000100101", -- i=212, alt=37, thresh=3.70908e-009, actual=7.2443e-012, err=0
        "0001010100000110111001110000000110", -- i=213, alt=6, thresh=3.01358e-009, actual=5.8859e-012, err=8.07794e-028
        "0110100001111011001111110000110011", -- i=214, alt=51, thresh=2.44611e-009, actual=4.77755e-012, err=8.07794e-028
        "0000101111110001010000010000001110", -- i=215, alt=14, thresh=1.98355e-009, actual=3.87412e-012, err=0
        "0011100111010111010010101000000101", -- i=216, alt=5, thresh=1.60689e-009, actual=3.13846e-012, err=4.03897e-028
        "0110011110101111011101100000101001", -- i=217, alt=41, thresh=1.30049e-009, actual=2.54001e-012, err=0
        "0110010110111111111011110000011000", -- i=218, alt=24, thresh=1.05148e-009, actual=2.05367e-012, err=0
        "0100100001011110101110000000000100", -- i=219, alt=4, thresh=8.4932e-010, actual=1.65883e-012, err=2.01948e-028
        "0101101001001011011000000000010011", -- i=220, alt=19, thresh=6.85358e-010, actual=1.33859e-012, err=0
        "0000010100000110011010001000011100", -- i=221, alt=28, thresh=5.52508e-010, actual=1.07912e-012, err=2.01948e-028
        "0010001111010101101110110000000011", -- i=222, alt=3, thresh=4.44975e-010, actual=8.69093e-013, err=0
        "0110010101110011001101111000100000", -- i=223, alt=32, thresh=3.58021e-010, actual=6.9926e-013, err=0
        "0100010010011010100100010000000010", -- i=224, alt=2, thresh=2.87778e-010, actual=5.62066e-013, err=0
        "0001101110001000000011101000101101", -- i=225, alt=45, thresh=2.3109e-010, actual=4.51348e-013, err=0
        "0100101110001101010110000000001101", -- i=226, alt=13, thresh=1.85388e-010, actual=3.62085e-013, err=0
        "0111110011000101101001001000000001", -- i=227, alt=1, thresh=1.48579e-010, actual=2.90193e-013, err=0
        "0010000110110110011101110000110010", -- i=228, alt=50, thresh=1.18962e-010, actual=2.32347e-013, err=0
        "0100111000101111010011000000100100", -- i=229, alt=36, thresh=9.51554e-011, actual=1.8585e-013, err=2.52435e-029
        "0010100111010000000100110000101000", -- i=230, alt=40, thresh=7.60389e-011, actual=1.48513e-013, err=2.52435e-029
        "0010000011110111010010100000010111", -- i=231, alt=23, thresh=6.07035e-011, actual=1.18561e-013, err=2.52435e-029
        "0001111000011101110101011000010010", -- i=232, alt=18, thresh=4.84135e-011, actual=9.45577e-014, err=1.26218e-029
        "0110101100111111011110100000001100", -- i=233, alt=12, thresh=3.85741e-011, actual=7.534e-014, err=0
        "0100110100110000110011101000011011", -- i=234, alt=27, thresh=3.07044e-011, actual=5.99695e-014, err=1.26218e-029
        "0010101100011010101000100000110001", -- i=235, alt=49, thresh=2.44163e-011, actual=4.76881e-014, err=6.31089e-030
        "0101010110011101110000100000101100", -- i=236, alt=44, thresh=1.93971e-011, actual=3.78849e-014, err=6.31089e-030
        "0110100101001001100010101000011111", -- i=237, alt=31, thresh=1.53946e-011, actual=3.00675e-014, err=6.31089e-030
        "0111111011010000001110000000100011", -- i=238, alt=35, thresh=1.2206e-011, actual=2.38399e-014, err=3.15544e-030
        "0000010111000011111011001000001011", -- i=239, alt=11, thresh=9.66845e-012, actual=1.88837e-014, err=0
        "0110100101011011010101100000100111", -- i=240, alt=39, thresh=7.65094e-012, actual=1.49433e-014, err=0
        "0011100111011111001101011000010110", -- i=241, alt=22, thresh=6.04852e-012, actual=1.18135e-014, err=0
        "0011100001100000111010000000010001", -- i=242, alt=17, thresh=4.77703e-012, actual=9.33014e-015, err=1.57772e-030
        "0111011100000001100111010000110000", -- i=243, alt=48, thresh=3.76915e-012, actual=7.36162e-015, err=0
        "0010101000011011000100101000001010", -- i=244, alt=10, thresh=2.97101e-012, actual=5.80275e-015, err=7.88861e-031
        "0011100011101110001011010000101011", -- i=245, alt=43, thresh=2.33959e-012, actual=4.56951e-015, err=7.88861e-031
        "0010111100010000110011011000011010", -- i=246, alt=26, thresh=1.84057e-012, actual=3.59486e-015, err=0
        "0001100110010100010011010000011110", -- i=247, alt=30, thresh=1.44657e-012, actual=2.82533e-015, err=0
        "0100101000101010010111101000100010", -- i=248, alt=34, thresh=1.1358e-012, actual=2.21836e-015, err=3.9443e-031
        "0011010111001001100110010000010000", -- i=249, alt=16, thresh=8.90925e-013, actual=1.74009e-015, err=1.97215e-031
        "0011101000101010010011000000001001", -- i=250, alt=9, thresh=6.98161e-013, actual=1.36359e-015, err=0
        "0111110001000000000101111000010101", -- i=251, alt=21, thresh=5.46569e-013, actual=1.06752e-015, err=0
        "0010110100011001101001100000100110", -- i=252, alt=38, thresh=4.27475e-013, actual=8.34912e-016, err=9.86076e-032
        "0100000101011101001110000000101111", -- i=253, alt=47, thresh=3.34004e-013, actual=6.52352e-016, err=0
        "0101100111100101110100010000001000", -- i=254, alt=8, thresh=2.60716e-013, actual=5.09212e-016, err=0
        "0000000011101011011010000000000000", -- i=255, alt=0, thresh=2.03311e-013, actual=3.97092e-016, err=0
        "0011000010100101110001001000101010", -- i=256, alt=42, thresh=1.5839e-013, actual=3.09356e-016, err=4.93038e-032
        "0000010100111101001010000000011001", -- i=257, alt=25, thresh=1.23274e-013, actual=2.4077e-016, err=0
        "0011100100100001101100001000001111", -- i=258, alt=15, thresh=9.58498e-014, actual=1.87207e-016, err=0
        "0011111000110010011101000000011101", -- i=259, alt=29, thresh=7.44537e-014, actual=1.45417e-016, err=2.46519e-032
        "0000000100011010101000110000000111", -- i=260, alt=7, thresh=5.77772e-014, actual=1.12846e-016, err=2.46519e-032
        "0101000000101110110000000000100001", -- i=261, alt=33, thresh=4.47922e-014, actual=8.74848e-017, err=1.2326e-032
        "0110000111101101111100011000010100", -- i=262, alt=20, thresh=3.46916e-014, actual=6.7757e-017, err=1.2326e-032
        "0011100010100011011110100000101110", -- i=263, alt=46, thresh=2.68424e-014, actual=5.24265e-017, err=0
        "0101101101111100010000000000100101", -- i=264, alt=37, thresh=2.07488e-014, actual=4.05251e-017, err=0
        "0011110001101110001010000000000110", -- i=265, alt=6, thresh=1.60229e-014, actual=3.12948e-017, err=0
        "0101100010101100010111110000001110", -- i=266, alt=14, thresh=1.23614e-014, actual=2.41433e-017, err=3.08149e-033
        "0111101010001000010100101000000101", -- i=267, alt=5, thresh=9.52721e-015, actual=1.86078e-017, err=0
        "0110000001101001010110111000101001", -- i=268, alt=41, thresh=7.33569e-015, actual=1.43275e-017, err=0
        "0110000100110011110010001000011000", -- i=269, alt=24, thresh=5.64276e-015, actual=1.1021e-017, err=1.54074e-033
        "0001111100101001111000010000000100", -- i=270, alt=4, thresh=4.33629e-015, actual=8.46932e-018, err=0
        "0001111100100000111000011000010011", -- i=271, alt=19, thresh=3.32905e-015, actual=6.50205e-018, err=0
        "0111100010110011100001100000011100", -- i=272, alt=28, thresh=2.55328e-015, actual=4.98687e-018, err=7.70372e-034
        "0100001011111101000110110000000011", -- i=273, alt=3, thresh=1.95637e-015, actual=3.82104e-018, err=7.70372e-034
        "0100011011111101000010001000100000", -- i=274, alt=32, thresh=1.49755e-015, actual=2.92489e-018, err=0
        "0101110110000011101111101000000010", -- i=275, alt=2, thresh=1.14521e-015, actual=2.23674e-018, err=0
        "0110110000010001110101100000101101", -- i=276, alt=45, thresh=8.74913e-016, actual=1.70881e-018, err=1.92593e-034
        "0111110110010010110001111000001101", -- i=277, alt=13, thresh=6.6776e-016, actual=1.30422e-018, err=1.92593e-034
        "0010110111000010110000100000000001", -- i=278, alt=1, thresh=5.09157e-016, actual=9.94447e-019, err=0
        "0010110111011000100110100000100100", -- i=279, alt=36, thresh=3.87845e-016, actual=7.57511e-019, err=0
        "0111001001000001100001011000101000", -- i=280, alt=40, thresh=2.95149e-016, actual=5.76463e-019, err=0
        "0110100100101010110011110000010111", -- i=281, alt=23, thresh=2.24388e-016, actual=4.38258e-019, err=0
        "0001000011011111000101111000010010", -- i=282, alt=18, thresh=1.70425e-016, actual=3.32861e-019, err=4.81482e-035
        "0000011100111011001101100000001100", -- i=283, alt=12, thresh=1.29313e-016, actual=2.52565e-019, err=0
        "0011011100111100101110111000011011", -- i=284, alt=27, thresh=9.80229e-017, actual=1.91451e-019, err=0
        "0001100110101110000010111000101100", -- i=285, alt=44, thresh=7.42315e-017, actual=1.44983e-019, err=0
        "0101001111101101110010001000011111", -- i=286, alt=31, thresh=5.61596e-017, actual=1.09687e-019, err=2.40741e-035
        "0001111101010100111000010000100011", -- i=287, alt=35, thresh=4.24459e-017, actual=8.29022e-020, err=1.20371e-035
        "0010001110010101011100110000001011", -- i=288, alt=11, thresh=3.20497e-017, actual=6.2597e-020, err=0
        "0111010001001001110010001000100111", -- i=289, alt=39, thresh=2.41761e-017, actual=4.7219e-020, err=6.01853e-036
        "0000010000100101100110000000010110", -- i=290, alt=22, thresh=1.8219e-017, actual=3.5584e-020, err=0
        "0111100000111101001100010000010001", -- i=291, alt=17, thresh=1.37164e-017, actual=2.67898e-020, err=0
        "0010111101101101011100110000001010", -- i=292, alt=10, thresh=1.03164e-017, actual=2.01493e-020, err=0
        "0100010101111011010101100000101011", -- i=293, alt=43, thresh=7.75166e-018, actual=1.514e-020, err=0
        "0101100011011101100101101000011010", -- i=294, alt=26, thresh=5.81883e-018, actual=1.13649e-020, err=1.50463e-036
        "0011100010101110001100000000011110", -- i=295, alt=30, thresh=4.36367e-018, actual=8.5228e-021, err=1.50463e-036
        "0011011001000101110010100000100010", -- i=296, alt=34, thresh=3.26922e-018, actual=6.3852e-021, err=7.52316e-037
        "0100011000110110000011110000010000", -- i=297, alt=16, thresh=2.44688e-018, actual=4.77906e-021, err=0
        "0000011011001100011110010000001001", -- i=298, alt=9, thresh=1.8296e-018, actual=3.57344e-021, err=7.52316e-037
        "0011001101110001101110001000010101", -- i=299, alt=21, thresh=1.36671e-018, actual=2.66935e-021, err=0
        "0011100000000010001000101000100110", -- i=300, alt=38, thresh=1.01993e-018, actual=1.99205e-021, err=0
        "0110011010101100110101111000001000", -- i=301, alt=8, thresh=7.60396e-019, actual=1.48515e-021, err=1.88079e-037
        "0110000110001001001111011000000000", -- i=302, alt=0, thresh=5.66351e-019, actual=1.10615e-021, err=0
        "0001110101111010100100000000101010", -- i=303, alt=42, thresh=4.21413e-019, actual=8.23071e-022, err=9.40395e-038
        "0011100101001110000001100000011001", -- i=304, alt=25, thresh=3.1326e-019, actual=6.11835e-022, err=9.40395e-038
        "0100110111010100011110100000001111", -- i=305, alt=15, thresh=2.32636e-019, actual=4.54368e-022, err=0
        "0010111010010001000011110000011101", -- i=306, alt=29, thresh=1.72594e-019, actual=3.37098e-022, err=4.70198e-038
        "0010100010100010000101001000000111", -- i=307, alt=7, thresh=1.27923e-019, actual=2.4985e-022, err=4.70198e-038
        "0111101111100010111011100000100001", -- i=308, alt=33, thresh=9.47217e-020, actual=1.85003e-022, err=2.35099e-038
        "0110100101101000011111001000010100", -- i=309, alt=20, thresh=7.00688e-020, actual=1.36853e-022, err=2.35099e-038
        "0011110001111010010001111000100101", -- i=310, alt=37, thresh=5.17816e-020, actual=1.01136e-022, err=0
        "0011010000011001001110101000000110", -- i=311, alt=6, thresh=3.82298e-020, actual=7.46675e-023, err=1.17549e-038
        "0100111001100010010010000000001110", -- i=312, alt=14, thresh=2.81971e-020, actual=5.50724e-023, err=1.17549e-038
        "0000001010010100111101011000000101", -- i=313, alt=5, thresh=2.07769e-020, actual=4.05799e-023, err=5.87747e-039
        "0110000111111101000111010000101001", -- i=314, alt=41, thresh=1.52945e-020, actual=2.9872e-023, err=0
        "0010000010011001111010111000011000", -- i=315, alt=24, thresh=1.12477e-020, actual=2.19681e-023, err=0
        "0011101101110111100110101000000100", -- i=316, alt=4, thresh=8.26357e-021, actual=1.61398e-023, err=2.93874e-039
        "0110111111100111001000101000010011", -- i=317, alt=19, thresh=6.06524e-021, actual=1.18462e-023, err=0
        "0101100011111010011111100000011100", -- i=318, alt=28, thresh=4.44737e-021, actual=8.68628e-024, err=1.46937e-039
        "0101001011100000110011110000000011", -- i=319, alt=3, thresh=3.25788e-021, actual=6.36304e-024, err=7.34684e-040
        "0000001100000110110001101000100000", -- i=320, alt=32, thresh=2.3842e-021, actual=4.65663e-024, err=7.34684e-040
        "0001111110100011110001011000000010", -- i=321, alt=2, thresh=1.74311e-021, actual=3.40451e-024, err=0
        "0010100010010001010000001000001101", -- i=322, alt=13, thresh=1.27316e-021, actual=2.48664e-024, err=3.67342e-040
        "0100110100000101111110010000000001", -- i=323, alt=1, thresh=9.29001e-022, actual=1.81445e-024, err=0
        "0010101000110000111000101000100100", -- i=324, alt=36, thresh=6.77213e-022, actual=1.32268e-024, err=0
        "0100000010011100111011111000101000", -- i=325, alt=40, thresh=4.93186e-022, actual=9.63253e-025, err=1.83671e-040
        "0000100010110100000001110000010111", -- i=326, alt=23, thresh=3.58815e-022, actual=7.00811e-025, err=0
        "0011100111011101011111111000010010", -- i=327, alt=18, thresh=2.608e-022, actual=5.09374e-025, err=9.18355e-041
        "0000010001101101111001001000001100", -- i=328, alt=12, thresh=1.89373e-022, actual=3.6987e-025, err=4.59177e-041
        "0001101011001101111100001000011011", -- i=329, alt=27, thresh=1.37375e-022, actual=2.6831e-025, err=4.59177e-041
        "0101111110111110100001110000011111", -- i=330, alt=31, thresh=9.95564e-023, actual=1.94446e-025, err=2.29589e-041
        "0001110111111110111101011000100011", -- i=331, alt=35, thresh=7.20789e-023, actual=1.40779e-025, err=0
        "0000110001111100001101111000001011", -- i=332, alt=11, thresh=5.21341e-023, actual=1.01824e-025, err=1.14794e-041
        "0101011001111100100110111000100111", -- i=333, alt=39, thresh=3.76714e-023, actual=7.3577e-026, err=0
        "0111100111000110111010011000010110", -- i=334, alt=22, thresh=2.71943e-023, actual=5.31138e-026, err=0
        "0111010111001011010000100000010001", -- i=335, alt=17, thresh=1.96118e-023, actual=3.83044e-026, err=5.73972e-042
        "0001000101101110011011110000001010", -- i=336, alt=10, thresh=1.41298e-023, actual=2.75972e-026, err=0
        "0000101011111100001010000000011010", -- i=337, alt=26, thresh=1.01701e-023, actual=1.98636e-026, err=0
        "0011000111100100011000011000011110", -- i=338, alt=30, thresh=7.31299e-024, actual=1.42832e-026, err=0
        "0101001011100111000100110000100010", -- i=339, alt=34, thresh=5.25338e-024, actual=1.02605e-026, err=0
        "0111100100010001011011010000010000", -- i=340, alt=16, thresh=3.77014e-024, actual=7.36356e-027, err=0
        "0011010000000010010111010000001001", -- i=341, alt=9, thresh=2.70304e-024, actual=5.27937e-027, err=7.17465e-043
        "0101010111111111000110110000010101", -- i=342, alt=21, thresh=1.93608e-024, actual=3.7814e-027, err=7.17465e-043
        "0001001010101001100100101000100110", -- i=343, alt=38, thresh=1.38538e-024, actual=2.70582e-027, err=0
        "0100011001101111111001010000001000", -- i=344, alt=8, thresh=9.90353e-025, actual=1.93428e-027, err=3.58732e-043
        "0100001101010001011110101000000000", -- i=345, alt=0, thresh=7.07273e-025, actual=1.38139e-027, err=1.79366e-043
        "0100100001001001100111011000011001", -- i=346, alt=25, thresh=5.04615e-025, actual=9.85576e-028, err=0
        "0111101000000111000100001000001111", -- i=347, alt=15, thresh=3.59673e-025, actual=7.02487e-028, err=8.96831e-044
        "0001011110011100110011100000011101", -- i=348, alt=29, thresh=2.56113e-025, actual=5.00221e-028, err=8.96831e-044
        "0011000101011100010100101000000111", -- i=349, alt=7, thresh=1.82193e-025, actual=3.55846e-028, err=4.48416e-044
        "0000010000010000011000100000100001", -- i=350, alt=33, thresh=1.29481e-025, actual=2.52893e-028, err=4.48416e-044
        "0010001100111110101101110000010100", -- i=351, alt=20, thresh=9.19301e-026, actual=1.79551e-028, err=0
        "0000011011100010011100101000100101", -- i=352, alt=37, thresh=6.52055e-026, actual=1.27354e-028, err=2.24208e-044
        "0001110111000011101100110000000110", -- i=353, alt=6, thresh=4.62047e-026, actual=9.02436e-029, err=1.12104e-044
        "0101010111111010010110111000001110", -- i=354, alt=14, thresh=3.27087e-026, actual=6.38843e-029, err=0
        "0100101011111010000111100000000101", -- i=355, alt=5, thresh=2.31322e-026, actual=4.51801e-029, err=5.60519e-045
        "0000010001001111001000010000011000", -- i=356, alt=24, thresh=1.63435e-026, actual=3.1921e-029, err=5.60519e-045
        "0111111110100010100010001000000100", -- i=357, alt=4, thresh=1.15359e-026, actual=2.2531e-029, err=2.8026e-045
        "0110001001011111100011001000010011", -- i=358, alt=19, thresh=8.13449e-027, actual=1.58877e-029, err=0
        "0110011100000111100111111000011100", -- i=359, alt=28, thresh=5.73041e-027, actual=1.11922e-029, err=0
        "0101001011111111010010110000000011", -- i=360, alt=3, thresh=4.0329e-027, actual=7.87676e-030, err=1.4013e-045
        "0000001001000011111011011000100000", -- i=361, alt=32, thresh=2.83546e-027, actual=5.53802e-030, err=0
        "0011101100000000101001001000000010", -- i=362, alt=2, thresh=1.99162e-027, actual=3.88988e-030, err=7.00649e-046
        "0000100010110110011111011000001101", -- i=363, alt=13, thresh=1.39754e-027, actual=2.72957e-030, err=3.50325e-046
        "0010011110101011000010011000000001", -- i=364, alt=1, thresh=9.79712e-028, actual=1.9135e-030, err=3.50325e-046
        "0110000001001001110001111000100100", -- i=365, alt=36, thresh=6.86132e-028, actual=1.3401e-030, err=0
        "0101001010110010000111110000010111", -- i=366, alt=23, thresh=4.80057e-028, actual=9.37611e-031, err=1.75162e-046
        "0011011111000001101101001000010010", -- i=367, alt=18, thresh=3.35547e-028, actual=6.55365e-031, err=0
        "0101101111011010011000101000001100", -- i=368, alt=12, thresh=2.34309e-028, actual=4.57635e-031, err=8.75812e-047
        "0110001100000110010100101000011011", -- i=369, alt=27, thresh=1.63456e-028, actual=3.1925e-031, err=4.37906e-047
        "0111100001010000011011000000011111", -- i=370, alt=31, thresh=1.13917e-028, actual=2.22494e-031, err=0
        "0000010111110011111001110000100011", -- i=371, alt=35, thresh=7.93143e-029, actual=1.54911e-031, err=0
        "0000001101011011010000100000001011", -- i=372, alt=11, thresh=5.51684e-029, actual=1.07751e-031, err=2.18953e-047
        "0110111010101111010001011000010110", -- i=373, alt=22, thresh=3.83358e-029, actual=7.48746e-032, err=1.09476e-047
        "0101011000001011001101001000010001", -- i=374, alt=17, thresh=2.6613e-029, actual=5.19786e-032, err=0
        "0100100110000111001001100000001010", -- i=375, alt=10, thresh=1.84569e-029, actual=3.60487e-032, err=0
        "0001101100110110011011000000011010", -- i=376, alt=26, thresh=1.27879e-029, actual=2.49764e-032, err=5.47382e-048
        "0001111000001011001000011000011110", -- i=377, alt=30, thresh=8.85151e-030, actual=1.72881e-032, err=2.73691e-048
        "0111110010101011000100100000100010", -- i=378, alt=34, thresh=6.12082e-030, actual=1.19547e-032, err=1.36846e-048
        "0100101000101011100101011000010000", -- i=379, alt=16, thresh=4.22841e-030, actual=8.25862e-033, err=0
        "0010111000001110000000111000001001", -- i=380, alt=9, thresh=2.91824e-030, actual=5.69969e-033, err=0
        "0111001011111011101111011000010101", -- i=381, alt=21, thresh=2.01206e-030, actual=3.9298e-033, err=0
        "0001101000001100001000000000001000", -- i=382, alt=8, thresh=1.38591e-030, actual=2.70685e-033, err=0
        "0001110001010010111011010000011001", -- i=383, alt=25, thresh=9.53685e-031, actual=1.86267e-033, err=0
        "0011010111101010101010111000001111", -- i=384, alt=15, thresh=6.55618e-031, actual=1.2805e-033, err=0
        "0011111000011001110000010000011101", -- i=385, alt=29, thresh=4.50269e-031, actual=8.79432e-034, err=0
        "0001000010101100100001111000000111", -- i=386, alt=7, thresh=3.08937e-031, actual=6.03392e-034, err=8.55285e-050
        "0011000011011101110011000000100001", -- i=387, alt=33, thresh=2.11759e-031, actual=4.13592e-034, err=8.55285e-050
        "0100000111110110111000010000010100", -- i=388, alt=20, thresh=1.45008e-031, actual=2.83218e-034, err=4.27642e-050
        "0001100111010101010010110000000110", -- i=389, alt=6, thresh=9.92007e-032, actual=1.93751e-034, err=4.27642e-050
        "0001100111110111101110100000001110", -- i=390, alt=14, thresh=6.77976e-032, actual=1.32417e-034, err=0
        "0000101001101001010100110000000101", -- i=391, alt=5, thresh=4.62902e-032, actual=9.04106e-035, err=0
        "0101001011000111100100100000011000", -- i=392, alt=24, thresh=3.15748e-032, actual=6.16695e-035, err=0
        "0000111111110011100100111000000100", -- i=393, alt=4, thresh=2.15162e-032, actual=4.20239e-035, err=5.34553e-051
        "0010000110010100011010001000010011", -- i=394, alt=19, thresh=1.46477e-032, actual=2.86087e-035, err=0
        "0111011001101111101011111000011100", -- i=395, alt=28, thresh=9.96199e-033, actual=1.9457e-035, err=2.67276e-051
        "0010101000001001001011010000000011", -- i=396, alt=3, thresh=6.76861e-033, actual=1.32199e-035, err=2.67276e-051
        "0010110010110000010000111000100000", -- i=397, alt=32, thresh=4.59439e-033, actual=8.97342e-036, err=1.33638e-051
        "0110010100101011000110010000000010", -- i=398, alt=2, thresh=3.11553e-033, actual=6.08503e-036, err=1.33638e-051
        "0001000111101001000111001000001101", -- i=399, alt=13, thresh=2.11063e-033, actual=4.12233e-036, err=0
        "0101101010110000001111000000000001", -- i=400, alt=1, thresh=1.42846e-033, actual=2.78996e-036, err=0
        "0100111011001010000110100000010111", -- i=401, alt=23, thresh=9.65828e-034, actual=1.88638e-036, err=0
        "0111101100010011101011010000010010", -- i=402, alt=18, thresh=6.52389e-034, actual=1.2742e-036, err=0
        "0111000111011011100101101000001100", -- i=403, alt=12, thresh=4.40239e-034, actual=8.59843e-037, err=0
        "0111001000100110000100100000011011", -- i=404, alt=27, thresh=2.96789e-034, actual=5.79665e-037, err=8.35239e-053
        "0110000111011010101100000000011111", -- i=405, alt=31, thresh=1.99885e-034, actual=3.90401e-037, err=0
        "0110101101100100110001110000001011", -- i=406, alt=11, thresh=1.3449e-034, actual=2.62676e-037, err=0
        "0011011110101010011011010000010110", -- i=407, alt=22, thresh=9.04014e-035, actual=1.76565e-037, err=0
        "0111011110100100111001000000010001", -- i=408, alt=17, thresh=6.07066e-035, actual=1.18568e-037, err=0
        "0111011100100001000100101000001010", -- i=409, alt=10, thresh=4.0726e-035, actual=7.9543e-038, err=0
        "0111100011101101001100111000011010", -- i=410, alt=26, thresh=2.7295e-035, actual=5.33106e-038, err=0
        "0111001010110001111100100000011110", -- i=411, alt=30, thresh=1.82756e-035, actual=3.56945e-038, err=5.22024e-054
        "0011010011111000100001100000010000", -- i=412, alt=16, thresh=1.22246e-035, actual=2.38761e-038, err=0
        "0011100110000100011001011000001001", -- i=413, alt=9, thresh=8.16907e-036, actual=1.59552e-038, err=0
        "0110100011011001100011101000010101", -- i=414, alt=21, thresh=5.45364e-036, actual=1.06516e-038, err=1.30506e-054
        "0101001010111011010111101000001000", -- i=415, alt=8, thresh=3.63728e-036, actual=7.10406e-039, err=1.30506e-054
        "0111110011111011101111000000011001", -- i=416, alt=25, thresh=2.42349e-036, actual=4.73339e-039, err=0
        "0001110101100111101110101000001111", -- i=417, alt=15, thresh=1.61318e-036, actual=3.15074e-039, err=6.5253e-055
        "0111111111111111111111111000011101", -- i=418, alt=29, thresh=0, actual=0, err=0
        "0111111111111111111111111000000111", -- i=419, alt=7, thresh=0, actual=0, err=0
        "0111111111111111111111111000010100", -- i=420, alt=20, thresh=0, actual=0, err=0
        "0111111111111111111111111000000110", -- i=421, alt=6, thresh=0, actual=0, err=0
        "0111111111111111111111111000001110", -- i=422, alt=14, thresh=0, actual=0, err=0
        "0111111111111111111111111000000101", -- i=423, alt=5, thresh=0, actual=0, err=0
        "0111111111111111111111111000011000", -- i=424, alt=24, thresh=0, actual=0, err=0
        "0111111111111111111111111000000100", -- i=425, alt=4, thresh=0, actual=0, err=0
        "0111111111111111111111111000010011", -- i=426, alt=19, thresh=0, actual=0, err=0
        "0111111111111111111111111000011100", -- i=427, alt=28, thresh=0, actual=0, err=0
        "0111111111111111111111111000000011", -- i=428, alt=3, thresh=0, actual=0, err=0
        "0111111111111111111111111000000010", -- i=429, alt=2, thresh=0, actual=0, err=0
        "0111111111111111111111111000001101", -- i=430, alt=13, thresh=0, actual=0, err=0
        "0111111111111111111111111000000001", -- i=431, alt=1, thresh=0, actual=0, err=0
        "0111111111111111111111111000010111", -- i=432, alt=23, thresh=0, actual=0, err=0
        "0111111111111111111111111000010010", -- i=433, alt=18, thresh=0, actual=0, err=0
        "0111111111111111111111111000001100", -- i=434, alt=12, thresh=0, actual=0, err=0
        "0111111111111111111111111000011011", -- i=435, alt=27, thresh=0, actual=0, err=0
        "0111111111111111111111111000001011", -- i=436, alt=11, thresh=0, actual=0, err=0
        "0111111111111111111111111000010110", -- i=437, alt=22, thresh=0, actual=0, err=0
        "0111111111111111111111111000010001", -- i=438, alt=17, thresh=0, actual=0, err=0
        "0111111111111111111111111000001010", -- i=439, alt=10, thresh=0, actual=0, err=0
        "0111111111111111111111111000011010", -- i=440, alt=26, thresh=0, actual=0, err=0
        "0111111111111111111111111000010000", -- i=441, alt=16, thresh=0, actual=0, err=0
        "0111111111111111111111111000001001", -- i=442, alt=9, thresh=0, actual=0, err=0
        "0111111111111111111111111000010101", -- i=443, alt=21, thresh=0, actual=0, err=0
        "0111111111111111111111111000001000", -- i=444, alt=8, thresh=0, actual=0, err=0
        "0111111111111111111111111000011001", -- i=445, alt=25, thresh=0, actual=0, err=0
        "0111111111111111111111111000001111", -- i=446, alt=15, thresh=0, actual=0, err=0
        "0111111111111111111111111000000111", -- i=447, alt=7, thresh=0, actual=0, err=0
        "0111111111111111111111111000010100", -- i=448, alt=20, thresh=0, actual=0, err=0
        "0111111111111111111111111000000110", -- i=449, alt=6, thresh=0, actual=0, err=0
        "0111111111111111111111111000001110", -- i=450, alt=14, thresh=0, actual=0, err=0
        "0111111111111111111111111000000101", -- i=451, alt=5, thresh=0, actual=0, err=0
        "0111111111111111111111111000011000", -- i=452, alt=24, thresh=0, actual=0, err=0
        "0111111111111111111111111000000100", -- i=453, alt=4, thresh=0, actual=0, err=0
        "0111111111111111111111111000010011", -- i=454, alt=19, thresh=0, actual=0, err=0
        "0111111111111111111111111000000011", -- i=455, alt=3, thresh=0, actual=0, err=0
        "0111111111111111111111111000000010", -- i=456, alt=2, thresh=0, actual=0, err=0
        "0111111111111111111111111000001101", -- i=457, alt=13, thresh=0, actual=0, err=0
        "0111111111111111111111111000000001", -- i=458, alt=1, thresh=0, actual=0, err=0
        "0111111111111111111111111000010111", -- i=459, alt=23, thresh=0, actual=0, err=0
        "0111111111111111111111111000010010", -- i=460, alt=18, thresh=0, actual=0, err=0
        "0111111111111111111111111000001100", -- i=461, alt=12, thresh=0, actual=0, err=0
        "0111111111111111111111111000001011", -- i=462, alt=11, thresh=0, actual=0, err=0
        "0111111111111111111111111000010110", -- i=463, alt=22, thresh=0, actual=0, err=0
        "0111111111111111111111111000010001", -- i=464, alt=17, thresh=0, actual=0, err=0
        "0111111111111111111111111000001010", -- i=465, alt=10, thresh=0, actual=0, err=0
        "0111111111111111111111111000010000", -- i=466, alt=16, thresh=0, actual=0, err=0
        "0111111111111111111111111000001001", -- i=467, alt=9, thresh=0, actual=0, err=0
        "0111111111111111111111111000010101", -- i=468, alt=21, thresh=0, actual=0, err=0
        "0111111111111111111111111000001000", -- i=469, alt=8, thresh=0, actual=0, err=0
        "0111111111111111111111111000001111", -- i=470, alt=15, thresh=0, actual=0, err=0
        "0111111111111111111111111000000111", -- i=471, alt=7, thresh=0, actual=0, err=0
        "0111111111111111111111111000010100", -- i=472, alt=20, thresh=0, actual=0, err=0
        "0111111111111111111111111000000110", -- i=473, alt=6, thresh=0, actual=0, err=0
        "0111111111111111111111111000001110", -- i=474, alt=14, thresh=0, actual=0, err=0
        "0111111111111111111111111000000101", -- i=475, alt=5, thresh=0, actual=0, err=0
        "0111111111111111111111111000000100", -- i=476, alt=4, thresh=0, actual=0, err=0
        "0111111111111111111111111000010011", -- i=477, alt=19, thresh=0, actual=0, err=0
        "0111111111111111111111111000000011", -- i=478, alt=3, thresh=0, actual=0, err=0
        "0111111111111111111111111000000010", -- i=479, alt=2, thresh=0, actual=0, err=0
        "0111111111111111111111111000001101", -- i=480, alt=13, thresh=0, actual=0, err=0
        "0111111111111111111111111000000001", -- i=481, alt=1, thresh=0, actual=0, err=0
        "0111111111111111111111111000010010", -- i=482, alt=18, thresh=0, actual=0, err=0
        "0111111111111111111111111000001100", -- i=483, alt=12, thresh=0, actual=0, err=0
        "0111111111111111111111111000001011", -- i=484, alt=11, thresh=0, actual=0, err=0
        "0111111111111111111111111000010001", -- i=485, alt=17, thresh=0, actual=0, err=0
        "0111111111111111111111111000001010", -- i=486, alt=10, thresh=0, actual=0, err=0
        "0111111111111111111111111000010000", -- i=487, alt=16, thresh=0, actual=0, err=0
        "0111111111111111111111111000001001", -- i=488, alt=9, thresh=0, actual=0, err=0
        "0111111111111111111111111000001000", -- i=489, alt=8, thresh=0, actual=0, err=0
        "0111111111111111111111111000001111", -- i=490, alt=15, thresh=0, actual=0, err=0
        "0111111111111111111111111000000111", -- i=491, alt=7, thresh=0, actual=0, err=0
        "0111111111111111111111111000000110", -- i=492, alt=6, thresh=0, actual=0, err=0
        "0111111111111111111111111000001110", -- i=493, alt=14, thresh=0, actual=0, err=0
        "0111111111111111111111111000000101", -- i=494, alt=5, thresh=0, actual=0, err=0
        "0111111111111111111111111000000100", -- i=495, alt=4, thresh=0, actual=0, err=0
        "0111111111111111111111111000000011", -- i=496, alt=3, thresh=0, actual=0, err=0
        "0111111111111111111111111000000010", -- i=497, alt=2, thresh=0, actual=0, err=0
        "0111111111111111111111111000001101", -- i=498, alt=13, thresh=0, actual=0, err=0
        "0111111111111111111111111000000001", -- i=499, alt=1, thresh=0, actual=0, err=0
        "0111111111111111111111111000001100", -- i=500, alt=12, thresh=0, actual=0, err=0
        "0111111111111111111111111000001011", -- i=501, alt=11, thresh=0, actual=0, err=0
        "0111111111111111111111111000001010", -- i=502, alt=10, thresh=0, actual=0, err=0
        "0111111111111111111111111000001001", -- i=503, alt=9, thresh=0, actual=0, err=0
        "0111111111111111111111111000001000", -- i=504, alt=8, thresh=0, actual=0, err=0
        "0111111111111111111111111000000111", -- i=505, alt=7, thresh=0, actual=0, err=0
        "0111111111111111111111111000000110", -- i=506, alt=6, thresh=0, actual=0, err=0
        "0111111111111111111111111000000101", -- i=507, alt=5, thresh=0, actual=0, err=0
        "0111111111111111111111111000000100", -- i=508, alt=4, thresh=0, actual=0, err=0
        "0111111111111111111111111000000011", -- i=509, alt=3, thresh=0, actual=0, err=0
        "0111111111111111111111111000000010", -- i=510, alt=2, thresh=0, actual=0, err=0
        "0111111111111111111111111000000001", -- i=511, alt=1, thresh=0, actual=0, err=0
        "0000000000010000100001110011111101", -- i=0, alt=60, thresh=0.983859, actual=0.012471, err=0
        "0000000011000000111011101101000101", -- i=1, alt=9, thresh=0.811589, actual=0.0249298, err=0
        "0000000010111011011000100000000010", -- i=2, alt=43, thresh=0.817009, actual=0.0248933, err=-3.46945e-018
        "0000000011000001110011100111100100", -- i=3, alt=21, thresh=0.810736, actual=0.0248326, err=0
        "0000000011001101001011111100110001", -- i=4, alt=68, thresh=0.799622, actual=0.0247478, err=0
        "0000000011001010110100110100001110", -- i=5, alt=59, thresh=0.801928, actual=0.0246392, err=0
        "0000000010111110011001001110111001", -- i=6, alt=30, thresh=0.814068, actual=0.0245071, err=0
        "0000000001011100110100000101111101", -- i=7, alt=22, thresh=0.909361, actual=0.024352, err=-3.46945e-018
        "0000000000010101000011011101010001", -- i=8, alt=25, thresh=0.979439, actual=0.0241741, err=3.46945e-018
        "0000000000000100110100110101010010", -- i=9, alt=25, thresh=0.995288, actual=0.0239742, err=0
        "0000000000010001010110110100000101", -- i=10, alt=53, thresh=0.98305, actual=0.0237526, err=0
        "0000000000000000111111100010101001", -- i=11, alt=34, thresh=0.99903, actual=0.0235102, err=0
        "0000000001001100110010110010100111", -- i=12, alt=16, thresh=0.925006, actual=0.0232474, err=0
        "0000000010111011110000100100111010", -- i=13, alt=26, thresh=0.816642, actual=0.0229652, err=3.46945e-018
        "0000000010110000100111010110011010", -- i=14, alt=48, thresh=0.827525, actual=0.0226642, err=0
        "0000000000000000000001010111111101", -- i=15, alt=60, thresh=0.999979, actual=0.0223454, err=0
        "0000000000000001111000010110110110", -- i=16, alt=53, thresh=0.998163, actual=0.0220095, err=0
        "0000000000011011110000101010010000", -- i=17, alt=67, thresh=0.97289, actual=0.0216574, err=0
        "0000000001001100010001001010101001", -- i=18, alt=61, thresh=0.925519, actual=0.0212902, err=0
        "0000000010110101111010100010001010", -- i=19, alt=8, thresh=0.822349, actual=0.0209088, err=0
        "0000000001111101010111000001000101", -- i=20, alt=21, thresh=0.877578, actual=0.0205141, err=0
        "0000000000001111111110100010001110", -- i=21, alt=30, thresh=0.984397, actual=0.0201073, err=0
        "0000000000000100011001010011000011", -- i=22, alt=35, thresh=0.995708, actual=0.0196892, err=0
        "0000000001110001001010111001100001", -- i=23, alt=71, thresh=0.889482, actual=0.019261, err=-3.46945e-018
        "0000000011100010000010011000001100", -- i=24, alt=8, thresh=0.779261, actual=0.0188238, err=0
        "0000000000000000010011111001111000", -- i=25, alt=61, thresh=0.999696, actual=0.0183785, err=-3.46945e-018
        "0000000000000010010011101111110010", -- i=26, alt=34, thresh=0.997746, actual=0.0179261, err=0
        "0000000000100111100010101101000101", -- i=27, alt=25, thresh=0.961385, actual=0.0174679, err=0
        "0000000010111111110000101111010010", -- i=28, alt=69, thresh=0.812733, actual=0.0170047, err=0
        "0000000000001111001100000001010111", -- i=29, alt=72, thresh=0.985168, actual=0.0165377, err=0
        "0000000000000001000010010100010101", -- i=30, alt=15, thresh=0.998988, actual=0.0160678, err=0
        "0000000000000011101111001101000101", -- i=31, alt=69, thresh=0.99635, actual=0.0155959, err=-1.73472e-018
        "0000000010110110000001100010111101", -- i=32, alt=0, thresh=0.822242, actual=0.0151232, err=1.73472e-018
        "0000000001011110100111111110000001", -- i=33, alt=9, thresh=0.907593, actual=0.0146504, err=1.73472e-018
        "0000000001011110100111111110000001", -- i=34, alt=34, thresh=NaN, actual=0.0141786, err=-7.45931e-017
        "0000000000000000111000110010101011", -- i=35, alt=60, thresh=0.999133, actual=0.0137085, err=1.73472e-018
        "0000000010111010011011100010110010", -- i=36, alt=10, thresh=0.817939, actual=0.0132411, err=-1.73472e-018
        "0000000010101011100111001100101111", -- i=37, alt=59, thresh=0.83241, actual=0.0127772, err=0
        "0000000000001110011001010100100010", -- i=38, alt=11, thresh=0.985942, actual=0.0123174, err=0
        "0000000000000010000001100001100001", -- i=39, alt=67, thresh=0.998024, actual=0.0118626, err=-1.73472e-018
        "0000000010000000010001101001100111", -- i=40, alt=52, thresh=0.874731, actual=0.0114135, err=0
        "0000000011011001110011100101110000", -- i=41, alt=47, thresh=0.787299, actual=0.0109706, err=0
        "0000000000010011010011110001011111", -- i=42, alt=39, thresh=0.981144, actual=0.0105346, err=-3.46945e-018
        "0000000000000101100000111100000011", -- i=43, alt=61, thresh=0.994615, actual=0.010106, err=-1.73472e-018
        "0000000000011101000110011100100100", -- i=44, alt=30, thresh=0.971581, actual=0.00968546, err=0
        "0000000010111111110100101000101010", -- i=45, alt=34, thresh=0.812673, actual=0.00927331, err=0
        "0000000010010001100001110010100000", -- i=46, alt=68, thresh=0.857883, actual=0.00887002, err=-1.73472e-018
        "0000000000001000000110111010011000", -- i=47, alt=39, thresh=0.992082, actual=0.00847599, err=0
        "0000000000011001111100100011011000", -- i=48, alt=35, thresh=0.974662, actual=0.00809155, err=1.73472e-018
        "0000000000100001110001111100110010", -- i=49, alt=11, thresh=0.967011, actual=0.00771701, err=0
        "0000000011000101010011111001101001", -- i=50, alt=38, thresh=0.807314, actual=0.00735261, err=8.67362e-019
        "0000000010110000110001010110000000", -- i=51, alt=42, thresh=0.827372, actual=0.00699858, err=0
        "0000000000001100111000101100100001", -- i=52, alt=54, thresh=0.987416, actual=0.00665508, err=-8.67362e-019
        "0000000000000000000000101101010000", -- i=53, alt=34, thresh=0.999989, actual=0.00632227, err=0
        "0000000000000000000111011100011000", -- i=54, alt=15, thresh=0.999886, actual=0.00600023, err=-8.67362e-019
        "0000000001000100111000001010101101", -- i=55, alt=54, thresh=0.932737, actual=0.00568903, err=0
        "0000000011000000110001010001101110", -- i=56, alt=16, thresh=0.811748, actual=0.00538871, err=0
        "0000000010111101010011000101000001", -- i=57, alt=60, thresh=0.815139, actual=0.00509925, err=0
        "0000000000110110111010001101011111", -- i=58, alt=34, thresh=0.946377, actual=0.00482063, err=8.67362e-019
        "0000000000100010100011110110001010", -- i=59, alt=69, thresh=0.96625, actual=0.00455279, err=8.67362e-019
        "0000000000000000000000010000010010", -- i=60, alt=34, thresh=0.999996, actual=0.00429562, err=0
        "0000000000000000000110010100100111", -- i=61, alt=67, thresh=0.999904, actual=0.00404902, err=0
        "0000000000100010011100110001110000", -- i=62, alt=53, thresh=0.966358, actual=0.00381285, err=0
        "0000000010000100000000101001010010", -- i=63, alt=38, thresh=0.871084, actual=0.00358695, err=-4.33681e-019
        "0000000010111111000010011101010001", -- i=64, alt=53, thresh=0.813439, actual=0.00337114, err=0
        "0000000011100101100000001000101010", -- i=65, alt=0, thresh=0.775877, actual=0.00316522, err=0
        "0000000010001010111101000000000001", -- i=66, alt=47, thresh=0.864304, actual=0.00296897, err=0
        "0000000000000000000010010100110110", -- i=67, alt=60, thresh=0.999965, actual=0.00278217, err=0
        "0000000000001001001010101000111010", -- i=68, alt=16, thresh=0.991049, actual=0.00260458, err=-4.33681e-019
        "0000000000000000010000101000001100", -- i=69, alt=54, thresh=0.999746, actual=0.00243594, err=-4.33681e-019
        "0000000000010001011000111010110001", -- i=70, alt=34, thresh=0.983018, actual=0.00227599, err=0
        "0000000000010111010101010111111101", -- i=71, alt=69, thresh=0.977213, actual=0.00212447, err=0
        "0000000000000000100001001011011001", -- i=72, alt=67, thresh=0.999494, actual=0.0019811, err=0
        "0000000000111000010111101111001000", -- i=73, alt=39, thresh=0.94495, actual=0.00184561, err=2.1684e-019
        "0000000001111011011011101100110100", -- i=74, alt=17, thresh=0.87946, actual=0.0017177, err=2.1684e-019
        "0000000010111010101010100110011101", -- i=75, alt=70, thresh=0.817709, actual=0.00159709, err=2.1684e-019
        "0000000011110110001110000001000110", -- i=76, alt=42, thresh=0.759552, actual=0.0014835, err=0
        "0000000100101110001111100001000110", -- i=77, alt=52, thresh=0.704841, actual=0.00137664, err=0
        "0000000101100010111000100111110010", -- i=78, alt=25, thresh=0.653433, actual=0.00127624, err=0
        "0000000110010100010010110001011010", -- i=79, alt=67, thresh=0.605182, actual=0.001182, err=2.1684e-019
        "0000000111000010100111010011010011", -- i=80, alt=15, thresh=0.559947, actual=0.00109365, err=2.1684e-019
        "0000000111101101111111011010000010", -- i=81, alt=29, thresh=0.517587, actual=0.00101091, err=0
        "0000001000101101001000001111111011", -- i=82, alt=58, thresh=0.477964, actual=0.000933524, err=0
        "0000001001111000111100100111011110", -- i=83, alt=7, thresh=0.440944, actual=0.000861218, err=1.0842e-019
        "0000001010111111101101001110010011", -- i=84, alt=33, thresh=0.406393, actual=0.000793737, err=0
        "0000001100000001101010111011111111", -- i=85, alt=20, thresh=0.374184, actual=0.000730828, err=1.0842e-019
        "0000001100111111000110001010010110", -- i=86, alt=66, thresh=0.344191, actual=0.000672249, err=0
        "0000001101111000001110110011110001", -- i=87, alt=46, thresh=0.316293, actual=0.00061776, err=0
        "0000001110101101010100010010000000", -- i=88, alt=37, thresh=0.290373, actual=0.000567134, err=1.0842e-019
        "0000001111011110100101011101000001", -- i=89, alt=6, thresh=0.266316, actual=0.000520148, err=0
        "0000010000011000100001010100100110", -- i=90, alt=51, thresh=0.244014, actual=0.000476589, err=0
        "0000010001101101000111011000011001", -- i=91, alt=14, thresh=0.223361, actual=0.000436251, err=5.42101e-020
        "0000010010111011010111100011001111", -- i=92, alt=57, thresh=0.204256, actual=0.000398937, err=5.42101e-020
        "0000010100000011101011001011101001", -- i=93, alt=5, thresh=0.186603, actual=0.000364459, err=5.42101e-020
        "0000010101000110011010100000111011", -- i=94, alt=41, thresh=0.170309, actual=0.000332635, err=0
        "0000010110000011111100101011100010", -- i=95, alt=65, thresh=0.155286, actual=0.000303293, err=0
        "0000010110111100100111101101101100", -- i=96, alt=24, thresh=0.14145, actual=0.00027627, err=0
        "0000010111110000110000100100010111", -- i=97, alt=4, thresh=0.128721, actual=0.000251408, err=5.42101e-020
        "0000011001000001010110010000110001", -- i=98, alt=19, thresh=0.117023, actual=0.00022856, err=0
        "0000011010011001010100011111101111", -- i=99, alt=28, thresh=0.106284, actual=0.000207586, err=0
        "0000011011101001111111011111100101", -- i=100, alt=3, thresh=0.0964365, actual=0.000188353, err=2.71051e-020
        "0000011100110011111000111011010101", -- i=101, alt=64, thresh=0.0874158, actual=0.000170734, err=0
        "0000011101110111100000100010111101", -- i=102, alt=32, thresh=0.0791616, actual=0.000154612, err=0
        "0000011110110101010100001111001101", -- i=103, alt=2, thresh=0.0716167, actual=0.000139876, err=2.71051e-020
        "0000011111101101110000000101110010", -- i=104, alt=45, thresh=0.0647276, actual=0.000126421, err=2.71051e-020
        "0000100001000010011100111011011000", -- i=105, alt=13, thresh=0.0584441, actual=0.000114149, err=1.35525e-020
        "0000100010100000010000000110111111", -- i=106, alt=56, thresh=0.052719, actual=0.000102967, err=0
        "0000100011110101100111111011110000", -- i=107, alt=1, thresh=0.0475083, actual=9.27897e-005, err=1.35525e-020
        "0000100101000011001111100100001001", -- i=108, alt=50, thresh=0.0427708, actual=8.35367e-005, err=0
        "0000100110001001101111010000110011", -- i=109, alt=36, thresh=0.0384681, actual=7.5133e-005, err=1.35525e-020
        "0000100111001001101100100001100000", -- i=110, alt=63, thresh=0.0345645, actual=6.75087e-005, err=1.35525e-020
        "0000101000000111010100011100000100", -- i=111, alt=40, thresh=0.0310266, actual=6.05989e-005, err=6.77626e-021
        "0000101001110000010001011101111000", -- i=112, alt=23, thresh=0.0278237, actual=5.43432e-005, err=0
        "0000101011001111001100001100011101", -- i=113, alt=18, thresh=0.024927, actual=4.86856e-005, err=0
        "0000101100100100111100001111011011", -- i=114, alt=12, thresh=0.0223101, actual=4.35745e-005, err=6.77626e-021
        "0000101101110010010101000010100001", -- i=115, alt=55, thresh=0.0199485, actual=3.89618e-005, err=0
        "0000101110111000000110000101100001", -- i=116, alt=27, thresh=0.0178194, actual=3.48034e-005, err=6.77626e-021
        "0000101111110110111011001011101101", -- i=117, alt=49, thresh=0.015902, actual=3.10585e-005, err=6.77626e-021
        "0000110001011110111001010101011010", -- i=118, alt=62, thresh=0.014177, actual=2.76895e-005, err=0
        "0000110011000100011111010001100100", -- i=119, alt=44, thresh=0.0126268, actual=2.46618e-005, err=3.38813e-021
        "0000110100011111101100010101001111", -- i=120, alt=31, thresh=0.0112352, actual=2.19437e-005, err=0
        "0000110101110001011111000000110101", -- i=121, alt=35, thresh=0.00998711, actual=1.95061e-005, err=3.38813e-021
        "0000110110111010110000100100110000", -- i=122, alt=11, thresh=0.00886903, actual=1.73223e-005, err=3.38813e-021
        "0000110111111100010101011001010001", -- i=123, alt=54, thresh=0.00786843, actual=1.5368e-005, err=0
        "0000111001101101111010101010010000", -- i=124, alt=61, thresh=0.0069739, actual=1.36209e-005, err=1.69407e-021
        "0000111011010110101000000101101100", -- i=125, alt=39, thresh=0.00617503, actual=1.20606e-005, err=1.69407e-021
        "0000111100110100000010101001111110", -- i=126, alt=22, thresh=0.00546233, actual=1.06686e-005, err=1.69407e-021
        "0000111110000111010010110010010101", -- i=127, alt=17, thresh=0.00482717, actual=9.42806e-006, err=1.69407e-021
        "0000111111010001011010010011111000", -- i=128, alt=48, thresh=0.0042617, actual=8.32362e-006, err=1.69407e-021
        "0001000000100110101001111110011111", -- i=129, alt=10, thresh=0.00375879, actual=7.34139e-006, err=8.47033e-022
        "0001000010011011110001111111111010", -- i=130, alt=43, thresh=0.00331199, actual=6.46873e-006, err=8.47033e-022
        "0001000100000011101110110011110001", -- i=131, alt=26, thresh=0.00291545, actual=5.69424e-006, err=8.47033e-022
        "0001000101011111111001001001010100", -- i=132, alt=60, thresh=0.00256389, actual=5.00759e-006, err=8.47033e-022
        "0001000110110001100001001010010110", -- i=133, alt=30, thresh=0.00225251, actual=4.39943e-006, err=0
        "0001000111111001101111001010101000", -- i=134, alt=53, thresh=0.00197702, actual=3.86136e-006, err=8.47033e-022
        "0001001001110011001000100111110110", -- i=135, alt=34, thresh=0.00173352, actual=3.38579e-006, err=4.23516e-022
        "0001001011100011110110011101010101", -- i=136, alt=16, thresh=0.00151853, actual=2.96589e-006, err=4.23516e-022
        "0001001101000111010001001111010110", -- i=137, alt=9, thresh=0.00132891, actual=2.59552e-006, err=0
        "0001001110011110110111100101101001", -- i=138, alt=21, thresh=0.00116183, actual=2.26919e-006, err=4.23516e-022
        "0001001111101011111110010110001001", -- i=139, alt=38, thresh=0.00101476, actual=1.98195e-006, err=4.23516e-022
        "0001010001011111100010111111011001", -- i=140, alt=59, thresh=0.000885442, actual=1.72938e-006, err=0
        "0001010011010110101010000000001111", -- i=141, alt=47, thresh=0.00077185, actual=1.50752e-006, err=2.11758e-022
        "0001010100111111001011001011010010", -- i=142, alt=8, thresh=0.000672174, actual=1.31284e-006, err=0
        "0001010110011010110010111000011000", -- i=143, alt=0, thresh=0.000584798, actual=1.14218e-006, err=2.11758e-022
        "0001010111101011000001101101011100", -- i=144, alt=42, thresh=0.000508283, actual=9.9274e-007, err=2.11758e-022
        "0001011001100010011011010011111011", -- i=145, alt=52, thresh=0.000441348, actual=8.62007e-007, err=0
        "0001011011011101000110010111001100", -- i=146, alt=25, thresh=0.000382853, actual=7.47759e-007, err=0
        "0001011101001000001100011001011000", -- i=147, alt=15, thresh=0.000331786, actual=6.4802e-007, err=1.05879e-022
        "0001011110100101100101111001110110", -- i=148, alt=29, thresh=0.00028725, actual=5.61036e-007, err=1.05879e-022
        "0001011111110110111101101001100000", -- i=149, alt=58, thresh=0.00024845, actual=4.85253e-007, err=0
        "0001100001111011100100001111011100", -- i=150, alt=7, thresh=0.00021468, actual=4.19297e-007, err=5.29396e-023
        "0001100011110110101101101101000101", -- i=151, alt=33, thresh=0.000185319, actual=3.61952e-007, err=5.29396e-023
        "0001100101100001101011001100111011", -- i=152, alt=20, thresh=0.000159818, actual=3.12144e-007, err=5.29396e-023
        "0001100110111110011110110101101101", -- i=153, alt=46, thresh=0.000137691, actual=2.68928e-007, err=5.29396e-023
        "0001101000011101110110011101110100", -- i=154, alt=37, thresh=0.000118512, actual=2.31468e-007, err=0
        "0001101010101001001010011110110101", -- i=155, alt=6, thresh=0.000101904, actual=1.99032e-007, err=2.64698e-023
        "0001101100100001101011000001010011", -- i=156, alt=51, thresh=8.75387e-005, actual=1.70974e-007, err=2.64698e-023
        "0001101110001001110011101111000001", -- i=157, alt=14, thresh=7.51247e-005, actual=1.46728e-007, err=2.64698e-023
        "0001101111100011101101000111110110", -- i=158, alt=57, thresh=6.44082e-005, actual=1.25797e-007, err=2.64698e-023
        "0001110001100010011101011111101000", -- i=159, alt=5, thresh=5.51664e-005, actual=1.07747e-007, err=1.32349e-023
        "0001110011101000000010011100000101", -- i=160, alt=41, thresh=4.72046e-005, actual=9.21965e-008, err=1.32349e-023
        "0001110101011010111111111011011011", -- i=161, alt=24, thresh=4.03524e-005, actual=7.88133e-008, err=1.32349e-023
        "0001110110111101110101100101011100", -- i=162, alt=4, thresh=3.44612e-005, actual=6.7307e-008, err=0
        "0001111000100101011101001100010001", -- i=163, alt=19, thresh=2.94013e-005, actual=5.74244e-008, err=0
        "0001111010110111001000011000101010", -- i=164, alt=28, thresh=2.50598e-005, actual=4.8945e-008, err=6.61744e-024
        "0001111100110011111111101100110100", -- i=165, alt=3, thresh=2.13386e-005, actual=4.1677e-008, err=6.61744e-024
        "0001111110011110111010011101100001", -- i=166, alt=32, thresh=1.81522e-005, actual=3.54535e-008, err=0
        "0001111111111010010111110011101111", -- i=167, alt=2, thresh=1.54265e-005, actual=3.01299e-008, err=6.61744e-024
        "0010000010010001000011011101111001", -- i=168, alt=45, thresh=1.30973e-005, actual=2.55807e-008, err=3.30872e-024
        "0010000100010110011111100000111000", -- i=169, alt=13, thresh=1.11089e-005, actual=2.16971e-008, err=0
        "0010000110001000010010100100011100", -- i=170, alt=56, thresh=9.41321e-006, actual=1.83852e-008, err=0
        "0010000111101001001111010111011101", -- i=171, alt=1, thresh=7.96854e-006, actual=1.55636e-008, err=0
        "0010001001110111100000011001001011", -- i=172, alt=50, thresh=6.739e-006, actual=1.31621e-008, err=0
        "0010001100000011110100001101110000", -- i=173, alt=36, thresh=5.69362e-006, actual=1.11203e-008, err=1.65436e-024
        "0010001101111010111111011001100110", -- i=174, alt=40, thresh=4.80569e-006, actual=9.38612e-009, err=1.65436e-024
        "0010001111100000000111001001111001", -- i=175, alt=23, thresh=4.05228e-006, actual=7.91462e-009, err=1.65436e-024
        "0010010001101011101001111100001010", -- i=176, alt=18, thresh=3.41365e-006, actual=6.66729e-009, err=8.27181e-025
        "0010010011111100110100101101101100", -- i=177, alt=12, thresh=2.87286e-006, actual=5.61105e-009, err=0
        "0010010101110111101000001100111101", -- i=178, alt=55, thresh=2.41537e-006, actual=4.71753e-009, err=8.27181e-025
        "0010010111011111011010001100101001", -- i=179, alt=27, thresh=2.02876e-006, actual=3.96242e-009, err=0
        "0010011001101110000011010001111001", -- i=180, alt=49, thresh=1.70236e-006, actual=3.32493e-009, err=0
        "0010011100000001110101110011010000", -- i=181, alt=44, thresh=1.42708e-006, actual=2.78727e-009, err=4.1359e-025
        "0010011101111110010110111111001011", -- i=182, alt=31, thresh=1.19515e-006, actual=2.33428e-009, err=4.1359e-025
        "0010011111100111001010100101100111", -- i=183, alt=35, thresh=9.99932e-007, actual=1.95299e-009, err=0
        "0010100001111110100101010001101100", -- i=184, alt=11, thresh=8.35785e-007, actual=1.63239e-009, err=0
        "0010100100010010101000100010111010", -- i=185, alt=54, thresh=6.97902e-007, actual=1.36309e-009, err=0
        "0010100110001110110111110000000100", -- i=186, alt=39, thresh=5.82197e-007, actual=1.1371e-009, err=2.06795e-025
        "0010100111110111000001010100101100", -- i=187, alt=22, thresh=4.852e-007, actual=9.47656e-010, err=2.06795e-025
        "0010101010011100011111000010011011", -- i=188, alt=17, thresh=4.03968e-007, actual=7.89e-010, err=0
        "0010101100101110011011011100101011", -- i=189, alt=48, thresh=3.36008e-007, actual=6.56265e-010, err=1.03398e-025
        "0010101110101000011010000001001100", -- i=190, alt=10, thresh=2.79207e-007, actual=5.45327e-010, err=0
        "0010110000011100100000001001101011", -- i=191, alt=43, thresh=2.31782e-007, actual=4.527e-010, err=0
        "0010110011000110011001101010001101", -- i=192, alt=26, thresh=1.92225e-007, actual=3.75439e-010, err=0
        "0010110101010011111110001110000100", -- i=193, alt=30, thresh=1.59263e-007, actual=3.1106e-010, err=0
        "0010110111001001110100100001110101", -- i=194, alt=53, thresh=1.31824e-007, actual=2.57469e-010, err=0
        "0010111001010111101001011001000110", -- i=195, alt=34, thresh=1.09006e-007, actual=2.12902e-010, err=0
        "0010111011111010011110110001001111", -- i=196, alt=16, thresh=9.00495e-008, actual=1.75878e-010, err=0
        "0010111110000001100111110010011110", -- i=197, alt=9, thresh=7.4317e-008, actual=1.4515e-010, err=0
        "0010111111110001101010101011011001", -- i=198, alt=21, thresh=6.12732e-008, actual=1.19674e-010, err=0
        "0011000010011100111100001011111100", -- i=199, alt=38, thresh=5.04695e-008, actual=9.85733e-011, err=1.29247e-026
        "0011000100110110100001001011011010", -- i=200, alt=47, thresh=4.15301e-008, actual=8.11135e-011, err=1.29247e-026
        "0011000110110101011101111010001100", -- i=201, alt=8, thresh=3.41407e-008, actual=6.6681e-011, err=0
        "0011001000111100100110010100000110", -- i=202, alt=0, thresh=2.80387e-008, actual=5.4763e-011, err=6.46235e-027
        "0011001011101001100011111101010010", -- i=203, alt=42, thresh=2.30048e-008, actual=4.49312e-011, err=6.46235e-027
        "0011001101111000000110110000111011", -- i=204, alt=52, thresh=1.88562e-008, actual=3.68285e-011, err=6.46235e-027
        "0011001111101101011101100110101010", -- i=205, alt=25, thresh=1.54407e-008, actual=3.01576e-011, err=6.46235e-027
        "0011010010011011111110001111001010", -- i=206, alt=15, thresh=1.26315e-008, actual=2.46708e-011, err=3.23117e-027
        "0011010100111010100101110101011001", -- i=207, alt=29, thresh=1.03233e-008, actual=2.01626e-011, err=3.23117e-027
        "0011010110111100110010100111111111", -- i=208, alt=7, thresh=8.4286e-009, actual=1.64621e-011, err=0
        "0011011001001111000111010001010111", -- i=209, alt=33, thresh=6.87495e-009, actual=1.34276e-011, err=0
        "0011011011111110000010011010000110", -- i=210, alt=20, thresh=5.60221e-009, actual=1.09418e-011, err=0
        "0011011110001101001100001111100000", -- i=211, alt=46, thresh=4.56063e-009, actual=8.90749e-012, err=1.61559e-027
        "0011100000000100011101001010000011", -- i=212, alt=37, thresh=3.70908e-009, actual=7.2443e-012, err=0
        "0011100011000011101000011111111110", -- i=213, alt=6, thresh=3.01358e-009, actual=5.8859e-012, err=8.07794e-028
        "0011100101011111100111101000101001", -- i=214, alt=51, thresh=2.44611e-009, actual=4.77755e-012, err=8.07794e-028
        "0011100111011110110001000000001011", -- i=215, alt=14, thresh=1.98355e-009, actual=3.87412e-012, err=0
        "0011101010001100100110011110111011", -- i=216, alt=5, thresh=1.60689e-009, actual=3.13846e-012, err=4.03897e-028
        "0011101100110101000011001011000011", -- i=217, alt=41, thresh=1.30049e-009, actual=2.54001e-012, err=0
        "0011101110111101111100010110010001", -- i=218, alt=24, thresh=1.05148e-009, actual=2.05367e-012, err=0
        "0011110001011010001010011011011110", -- i=219, alt=4, thresh=8.4932e-010, actual=1.65883e-012, err=2.01948e-028
        "0011110100001110011100001111100000", -- i=220, alt=19, thresh=6.85358e-010, actual=1.33859e-012, err=0
        "0011110110100000100000101011011011", -- i=221, alt=28, thresh=5.52508e-010, actual=1.07912e-012, err=2.01948e-028
        "0011111000101101011111010001000100", -- i=222, alt=3, thresh=4.44975e-010, actual=8.69093e-013, err=0
        "0011111011101100101100111110011010", -- i=223, alt=32, thresh=3.58021e-010, actual=6.9926e-013, err=0
        "0011111110000111001010110111101000", -- i=224, alt=2, thresh=2.87778e-010, actual=5.62066e-013, err=0
        "0100000000000111101001111010010101", -- i=225, alt=45, thresh=2.3109e-010, actual=4.51348e-013, err=0
        "0100000011010000101001111111000110", -- i=226, alt=13, thresh=1.85388e-010, actual=3.62085e-013, err=0
        "0100000101110010100010110101100111", -- i=227, alt=1, thresh=1.48579e-010, actual=2.90193e-013, err=0
        "0100000111110100110011010000011110", -- i=228, alt=50, thresh=1.18962e-010, actual=2.32347e-013, err=0
        "0100001010111011000000001111101111", -- i=229, alt=36, thresh=9.51554e-011, actual=1.8585e-013, err=2.52435e-029
        "0100001101100011001001111010011110", -- i=230, alt=40, thresh=7.60389e-011, actual=1.48513e-013, err=2.52435e-029
        "0100001111101010000010111111011100", -- i=231, alt=23, thresh=6.07035e-011, actual=1.18561e-013, err=2.52435e-029
        "0100010010101100010011001101101001", -- i=232, alt=18, thresh=4.84135e-011, actual=9.45577e-014, err=1.26218e-029
        "0100010101011001011001011100001010", -- i=233, alt=12, thresh=3.85741e-011, actual=7.534e-014, err=0
        "0100010111100011110101111101000110", -- i=234, alt=27, thresh=3.07044e-011, actual=5.99695e-014, err=1.26218e-029
        "0100011010100100111011010100110000", -- i=235, alt=49, thresh=2.44163e-011, actual=4.76881e-014, err=6.31089e-030
        "0100011101010101100001101100010000", -- i=236, alt=44, thresh=1.93971e-011, actual=3.78849e-014, err=6.31089e-030
        "0100011111100010010110100001100101", -- i=237, alt=31, thresh=1.53946e-011, actual=3.00675e-014, err=6.31089e-030
        "0100100010100101000100111100001011", -- i=238, alt=35, thresh=1.2206e-011, actual=2.38399e-014, err=3.15544e-030
        "0100100101010111101001001010110000", -- i=239, alt=11, thresh=9.66845e-012, actual=1.88837e-014, err=0
        "0100100111100101100111001101010010", -- i=240, alt=39, thresh=7.65094e-012, actual=1.49433e-014, err=0
        "0100101010101100101111110011110001", -- i=241, alt=22, thresh=6.04852e-012, actual=1.18135e-014, err=0
        "0100101101011111101100010011111101", -- i=242, alt=17, thresh=4.77703e-012, actual=9.33014e-015, err=1.57772e-030
        "0100101111101101100010100001110110", -- i=243, alt=48, thresh=3.76915e-012, actual=7.36162e-015, err=0
        "0100110010111011101111000100110001", -- i=244, alt=10, thresh=2.97101e-012, actual=5.80275e-015, err=7.88861e-031
        "0100110101101101011101101010011101", -- i=245, alt=43, thresh=2.33959e-012, actual=4.56951e-015, err=7.88861e-031
        "0100110111111001111011010001011101", -- i=246, alt=26, thresh=1.84057e-012, actual=3.59486e-015, err=0
        "0100111011010001101001110101101011", -- i=247, alt=30, thresh=1.44657e-012, actual=2.82533e-015, err=0
        "0100111110000000100110011100011110", -- i=248, alt=34, thresh=1.1358e-012, actual=2.21836e-015, err=3.9443e-031
        "0101000000010100111010000110110101", -- i=249, alt=16, thresh=8.90925e-013, actual=1.74009e-015, err=1.97215e-031
        "0101000011101101111100001110111100", -- i=250, alt=9, thresh=6.98161e-013, actual=1.36359e-015, err=0
        "0101000110011000100111100010011111", -- i=251, alt=21, thresh=5.46569e-013, actual=1.06752e-015, err=0
        "0101001000111101011010010111111001", -- i=252, alt=38, thresh=4.27475e-013, actual=8.34912e-016, err=9.86076e-032
        "0101001100001111111000111100100001", -- i=253, alt=47, thresh=3.34004e-013, actual=6.52352e-016, err=0
        "0101001110110100111010110011010100", -- i=254, alt=8, thresh=2.60716e-013, actual=5.09212e-016, err=0
        "0101010001101100010111100111011011", -- i=255, alt=0, thresh=2.03311e-013, actual=3.97092e-016, err=0
        "0101010100110110101011000110010111", -- i=256, alt=42, thresh=1.5839e-013, actual=3.09356e-016, err=4.93038e-032
        "0101010111010100110100101000100111", -- i=257, alt=25, thresh=1.23274e-013, actual=2.4077e-016, err=0
        "0101011010100000101010010101111110", -- i=258, alt=15, thresh=9.58498e-014, actual=1.87207e-016, err=0
        "0101011101100001011000011000111110", -- i=259, alt=29, thresh=7.44537e-014, actual=1.45417e-016, err=2.46519e-032
        "0101011111110111100101101110001010", -- i=260, alt=7, thresh=5.77772e-014, actual=1.12846e-016, err=2.46519e-032
        "0101100011011001000110000111100000", -- i=261, alt=33, thresh=4.47922e-014, actual=8.74848e-017, err=1.2326e-032
        "0101100110001111000011010110010011", -- i=262, alt=20, thresh=3.46916e-014, actual=6.7757e-017, err=1.2326e-032
        "0101101000111000111001101011011100", -- i=263, alt=46, thresh=2.68424e-014, actual=5.24265e-017, err=0
        "0101101100010100011100011011011100", -- i=264, alt=37, thresh=2.07488e-014, actual=4.05251e-017, err=0
        "0101101110111110101101100111001100", -- i=265, alt=6, thresh=1.60229e-014, actual=3.12948e-017, err=0
        "0101110010000101010001010010100010", -- i=266, alt=14, thresh=1.23614e-014, actual=2.41433e-017, err=3.08149e-033
        "0101110101010001011111011111001000", -- i=267, alt=5, thresh=9.52721e-015, actual=1.86078e-017, err=0
        "0101110111101111011010000101111010", -- i=268, alt=41, thresh=7.33569e-015, actual=1.43275e-017, err=0
        "0101111011010010110010101011111000", -- i=269, alt=24, thresh=5.64276e-015, actual=1.1021e-017, err=1.54074e-033
        "0101111110001111000100110010000001", -- i=270, alt=4, thresh=4.33629e-015, actual=8.46932e-018, err=0
        "0110000001000000011101110110110010", -- i=271, alt=19, thresh=3.32905e-015, actual=6.50205e-018, err=0
        "0110000100100000000100010101110000", -- i=272, alt=28, thresh=2.55328e-015, actual=4.98687e-018, err=7.70372e-034
        "0110000111001100000111010100010001", -- i=273, alt=3, thresh=1.95637e-015, actual=3.82104e-018, err=7.70372e-034
        "0110001010100000101110010011010110", -- i=274, alt=32, thresh=1.49755e-015, actual=2.92489e-018, err=0
        "0110001101101011110101010000001101", -- i=275, alt=2, thresh=1.14521e-015, actual=2.23674e-018, err=0
        "0110010000001111010010110101001100", -- i=276, alt=45, thresh=8.74913e-016, actual=1.70881e-018, err=1.92593e-034
        "0110010011111110001000000000000110", -- i=277, alt=13, thresh=6.6776e-016, actual=1.30422e-018, err=1.92593e-034
        "0110010110110100111110110101110000", -- i=278, alt=1, thresh=5.09157e-016, actual=9.94447e-019, err=0
        "0110011010000001101100000111011000", -- i=279, alt=36, thresh=3.87845e-016, actual=7.57511e-019, err=0
        "0110011101010111011011101101001000", -- i=280, alt=40, thresh=2.95149e-016, actual=5.76463e-019, err=0
        "0110011111111010100110001100100101", -- i=281, alt=23, thresh=2.24388e-016, actual=4.38258e-019, err=0
        "0110100011101110000011011100010001", -- i=282, alt=18, thresh=1.70425e-016, actual=3.32861e-019, err=4.81482e-035
        "0110100110101011101001100000111111", -- i=283, alt=12, thresh=1.29313e-016, actual=2.52565e-019, err=0
        "0110101001110111111001100000101000", -- i=284, alt=27, thresh=9.80229e-017, actual=1.91451e-019, err=0
        "0110101101010011010101011110110011", -- i=285, alt=44, thresh=7.42315e-017, actual=1.44983e-019, err=0
        "0110101111111010000001001101011110", -- i=286, alt=31, thresh=5.61596e-017, actual=1.09687e-019, err=2.40741e-035
        "0110110011110001000000101100110111", -- i=287, alt=35, thresh=4.24459e-017, actual=8.29022e-020, err=1.20371e-035
        "0110110110110000110010011100100000", -- i=288, alt=11, thresh=3.20497e-017, actual=6.2597e-020, err=0
        "0110111010000100000011110001111101", -- i=289, alt=39, thresh=2.41761e-017, actual=4.7219e-020, err=6.01853e-036
        "0110111101011111110101100011101011", -- i=290, alt=22, thresh=1.8219e-017, actual=3.5584e-020, err=0
        "0111000000001011111010010001010001", -- i=291, alt=17, thresh=1.37164e-017, actual=2.67898e-020, err=0
        "0111000100000110110010000101000101", -- i=292, alt=10, thresh=1.03164e-017, actual=2.01493e-020, err=0
        "0111000111000100000001110101101011", -- i=293, alt=43, thresh=7.75166e-018, actual=1.514e-020, err=0
        "0111001010100101010010101110000000", -- i=294, alt=26, thresh=5.81883e-018, actual=1.13649e-020, err=1.50463e-036
        "0111001101111100000010010001011001", -- i=295, alt=30, thresh=4.36367e-018, actual=8.5228e-021, err=1.50463e-036
        "0111010000111011000110001000011001", -- i=296, alt=34, thresh=3.26922e-018, actual=6.3852e-021, err=7.52316e-037
        "0111010100101101110011110001100111", -- i=297, alt=16, thresh=2.44688e-018, actual=4.77906e-021, err=0
        "0111010111100011111111110110110010", -- i=298, alt=9, thresh=1.8296e-018, actual=3.57344e-021, err=7.52316e-037
        "0111011011011001001111010100101100", -- i=299, alt=21, thresh=1.36671e-018, actual=2.66935e-021, err=0
        "0111011110100101111100001100100000", -- i=300, alt=38, thresh=1.01993e-018, actual=1.99205e-021, err=0
        "0111100001111110010010000101001000", -- i=301, alt=8, thresh=7.60396e-019, actual=1.48515e-021, err=1.88079e-037
        "0111100101100011010111101101000010", -- i=302, alt=0, thresh=5.66351e-019, actual=1.10615e-021, err=0
        "0111101000011100111101111011111110", -- i=303, alt=42, thresh=4.21413e-019, actual=8.23071e-022, err=9.40395e-038
        "0111101100011100010101100001100011", -- i=304, alt=25, thresh=3.1326e-019, actual=6.11835e-022, err=9.40395e-038
        "0111101111011010101101000000011001", -- i=305, alt=15, thresh=2.32636e-019, actual=4.54368e-022, err=0
        "0111110011010000111100101010010010", -- i=306, alt=29, thresh=1.72594e-019, actual=3.37098e-022, err=4.70198e-038
        "0111110110100011111001100011010001", -- i=307, alt=7, thresh=1.27923e-019, actual=2.4985e-022, err=4.70198e-038
        "0111111010000001011000010001011011", -- i=308, alt=33, thresh=9.47217e-020, actual=1.85003e-022, err=2.35099e-038
        "0111111101101010001110000001111000", -- i=309, alt=20, thresh=7.00688e-020, actual=1.36853e-022, err=2.35099e-038
        "1000000000101101110111111010100001", -- i=310, alt=37, thresh=5.17816e-020, actual=1.01136e-022, err=0
        "1000000100101101110111000010110100", -- i=311, alt=6, thresh=3.82298e-020, actual=7.46675e-023, err=1.17549e-038
        "1000000111101011010111110110110001", -- i=312, alt=14, thresh=2.81971e-020, actual=5.50724e-023, err=1.17549e-038
        "1000001011101111000100011110001000", -- i=313, alt=5, thresh=2.07769e-020, actual=4.05799e-023, err=5.87747e-039
        "1000001110111110001100001110101000", -- i=314, alt=41, thresh=1.52945e-020, actual=2.9872e-023, err=0
        "1000010010101110001001011111111001", -- i=315, alt=24, thresh=1.12477e-020, actual=2.19681e-023, err=0
        "1000010110001111100111110011111110", -- i=316, alt=4, thresh=8.26357e-021, actual=1.61398e-023, err=2.93874e-039
        "1000011001101011011100100110101011", -- i=317, alt=19, thresh=6.06524e-021, actual=1.18462e-023, err=0
        "1000011101011111111011101001000010", -- i=318, alt=28, thresh=4.44737e-021, actual=8.68628e-024, err=1.46937e-039
        "1000100000100111010111011101100100", -- i=319, alt=3, thresh=3.25788e-021, actual=6.36304e-024, err=7.34684e-040
        "1000100100101111011010111101011000", -- i=320, alt=32, thresh=2.3842e-021, actual=4.65663e-024, err=7.34684e-040
        "1000100111110001001011011000110010", -- i=321, alt=2, thresh=1.74311e-021, actual=3.40451e-024, err=0
        "1000101011111110011011000100101010", -- i=322, alt=13, thresh=1.27316e-021, actual=2.48664e-024, err=3.67342e-040
        "1000101111001110011101000001001010", -- i=323, alt=1, thresh=9.29001e-022, actual=1.81445e-024, err=0
        "1000110011001101010011001010001111", -- i=324, alt=36, thresh=6.77213e-022, actual=1.32268e-024, err=0
        "1000110110101011110001100111000100", -- i=325, alt=40, thresh=4.93186e-022, actual=9.63253e-025, err=1.83671e-040
        "1000111010011100011100000001010101", -- i=326, alt=23, thresh=3.58815e-022, actual=7.00811e-025, err=0
        "1000111110001001011011001100101011", -- i=327, alt=18, thresh=2.608e-022, actual=5.09374e-025, err=9.18355e-041
        "1001000001101100001111110010001000", -- i=328, alt=12, thresh=1.89373e-022, actual=3.6987e-025, err=4.59177e-041
        "1001000101100111101100101000110011", -- i=329, alt=27, thresh=1.37375e-022, actual=2.6831e-025, err=4.59177e-041
        "1001001000111101001001100100000001", -- i=330, alt=31, thresh=9.95564e-023, actual=1.94446e-025, err=2.29589e-041
        "1001001101000110111001010110100011", -- i=331, alt=35, thresh=7.20789e-023, actual=1.40779e-025, err=0
        "1001010000001111100101000101010110", -- i=332, alt=11, thresh=5.21341e-023, actual=1.01824e-025, err=1.14794e-041
        "1001010100100111010101000011011001", -- i=333, alt=39, thresh=3.76714e-023, actual=7.3577e-026, err=0
        "1001010111110001111111001000011101", -- i=334, alt=22, thresh=2.71943e-023, actual=5.31138e-026, err=0
        "1001011100001001010011011011111011", -- i=335, alt=17, thresh=1.96118e-023, actual=3.83044e-026, err=5.73972e-042
        "1001011111011101011000011001001001", -- i=336, alt=10, thresh=1.41298e-023, actual=2.75972e-026, err=0
        "1001100011101101000111110111101110", -- i=337, alt=26, thresh=1.01701e-023, actual=1.98636e-026, err=0
        "1001100111001010001011110100010100", -- i=338, alt=30, thresh=7.31299e-024, actual=1.42832e-026, err=0
        "1001101011010011000101000100101101", -- i=339, alt=34, thresh=5.25338e-024, actual=1.02605e-026, err=0
        "1001101110111000100110010100111001", -- i=340, alt=16, thresh=3.77014e-024, actual=7.36356e-027, err=0
        "1001110010111011011100110010101101", -- i=341, alt=9, thresh=2.70304e-024, actual=5.27937e-027, err=7.17465e-043
        "1001110110101000110100000010101100", -- i=342, alt=21, thresh=1.93608e-024, actual=3.7814e-027, err=7.17465e-043
        "1001111010100110011111011111010010", -- i=343, alt=38, thresh=1.38538e-024, actual=2.70582e-027, err=0
        "1001111110011011000000000100100000", -- i=344, alt=8, thresh=9.90353e-025, actual=1.93428e-027, err=3.58732e-043
        "1010000010010100011100000010101111", -- i=345, alt=0, thresh=7.07273e-025, actual=1.38139e-027, err=1.79366e-043
        "1010000110001111010100010011001011", -- i=346, alt=25, thresh=5.04615e-025, actual=9.85576e-028, err=0
        "1010001010000101011111011110100011", -- i=347, alt=15, thresh=3.59673e-025, actual=7.02487e-028, err=8.96831e-044
        "1010001110000101111001001101110100", -- i=348, alt=29, thresh=2.56113e-025, actual=5.00221e-028, err=8.96831e-044
        "1010010001111001110100101101110000", -- i=349, alt=7, thresh=1.82193e-025, actual=3.55846e-028, err=4.48416e-044
        "1010010101111110110101101111100001", -- i=350, alt=33, thresh=1.29481e-025, actual=2.52893e-028, err=4.48416e-044
        "1010011001110001100100010111100110", -- i=351, alt=20, thresh=9.19301e-026, actual=1.79551e-028, err=0
        "1010011101111010001111000110111011", -- i=352, alt=37, thresh=6.52055e-026, actual=1.27354e-028, err=2.24208e-044
        "1010100001101100110100100101000010", -- i=353, alt=6, thresh=4.62047e-026, actual=9.02436e-029, err=1.12104e-044
        "1010100101111000001000101111110000", -- i=354, alt=14, thresh=3.27087e-026, actual=6.38843e-029, err=0
        "1010101001101011101000111001000101", -- i=355, alt=5, thresh=2.31322e-026, actual=4.51801e-029, err=5.60519e-045
        "1010101101111000100100001110100101", -- i=356, alt=24, thresh=1.63435e-026, actual=3.1921e-029, err=5.60519e-045
        "1010110001101110000010001100011011", -- i=357, alt=4, thresh=1.15359e-026, actual=2.2531e-029, err=2.8026e-045
        "1010110101111011100001001110110010", -- i=358, alt=19, thresh=8.13449e-027, actual=1.58877e-029, err=0
        "1010111001110011111110101100010100", -- i=359, alt=28, thresh=5.73041e-027, actual=1.11922e-029, err=0
        "1010111110000000111101100011000101", -- i=360, alt=3, thresh=4.0329e-027, actual=7.87676e-030, err=1.4013e-045
        "1011000001111101011001111100110010", -- i=361, alt=32, thresh=2.83546e-027, actual=5.53802e-030, err=0
        "1011000110001000110101001000001010", -- i=362, alt=2, thresh=1.99162e-027, actual=3.88988e-030, err=7.00649e-046
        "1011001010001010001100111110001001", -- i=363, alt=13, thresh=1.39754e-027, actual=2.72957e-030, err=3.50325e-046
        "1011001110010011000010001001110000", -- i=364, alt=1, thresh=9.79712e-028, actual=1.9135e-030, err=3.50325e-046
        "1011010010011010001110010101101011", -- i=365, alt=36, thresh=6.86132e-028, actual=1.3401e-030, err=0
        "1011010110011111011101001001110010", -- i=366, alt=23, thresh=4.80057e-028, actual=9.37611e-031, err=1.75162e-046
        "1011011010101101010010011001001010", -- i=367, alt=18, thresh=3.35547e-028, actual=6.55365e-031, err=0
        "1011011110101101111101001001011111", -- i=368, alt=12, thresh=2.34309e-028, actual=4.57635e-031, err=8.75812e-047
        "1011100011000011001011011100111011", -- i=369, alt=27, thresh=1.63456e-028, actual=3.1925e-031, err=4.37906e-047
        "1011100110111110010111110100001011", -- i=370, alt=31, thresh=1.13917e-028, actual=2.22494e-031, err=0
        "1011101011011011101010000100010010", -- i=371, alt=35, thresh=7.93143e-029, actual=1.54911e-031, err=0
        "1011101111010000100001101011100000", -- i=372, alt=11, thresh=5.51684e-029, actual=1.07751e-031, err=2.18953e-047
        "1011110011110110011101010011100010", -- i=373, alt=22, thresh=3.83358e-029, actual=7.48746e-032, err=1.09476e-047
        "1011110111100100001110010100101101", -- i=374, alt=17, thresh=2.6613e-029, actual=5.19786e-032, err=0
        "1011111100010011010011000011100011", -- i=375, alt=10, thresh=1.84569e-029, actual=3.60487e-032, err=0
        "1011111111111001010000100110110101", -- i=376, alt=26, thresh=1.27879e-029, actual=2.49764e-032, err=5.47382e-048
        "1100000100110001111000010101111011", -- i=377, alt=30, thresh=8.85151e-030, actual=1.72881e-032, err=2.73691e-048
        "1100001000011110110101110010001011", -- i=378, alt=34, thresh=6.12082e-030, actual=1.19547e-032, err=1.36846e-048
        "1100001101010001111001101001101010", -- i=379, alt=16, thresh=4.22841e-030, actual=8.25862e-033, err=0
        "1100010001001100111110100011000110", -- i=380, alt=9, thresh=2.91824e-030, actual=5.69969e-033, err=0
        "1100010101110011000011001111101010", -- i=381, alt=21, thresh=2.01206e-030, actual=3.9298e-033, err=0
        "1100011001111100011111100110101111", -- i=382, alt=8, thresh=1.38591e-030, actual=2.70685e-033, err=0
        "1100011110010101000001011110100110", -- i=383, alt=25, thresh=9.53685e-031, actual=1.86267e-033, err=0
        "1100100010101100111101011001001000", -- i=384, alt=15, thresh=6.55618e-031, actual=1.2805e-033, err=0
        "1100100110110111100001000101101101", -- i=385, alt=29, thresh=4.50269e-031, actual=8.79432e-034, err=0
        "1100101011011101111101000101101110", -- i=386, alt=7, thresh=3.08937e-031, actual=6.03392e-034, err=8.55285e-050
        "1100101111011010001111011110010100", -- i=387, alt=33, thresh=2.11759e-031, actual=4.13592e-034, err=8.55285e-050
        "1100110100001111000100111110110101", -- i=388, alt=20, thresh=1.45008e-031, actual=2.83218e-034, err=4.27642e-050
        "1100110111111100111010111011011110", -- i=389, alt=6, thresh=9.92007e-032, actual=1.93751e-034, err=4.27642e-050
        "1100111100111111111100110010100010", -- i=390, alt=14, thresh=6.77976e-032, actual=1.32417e-034, err=0
        "1101000000111110100101101111010110", -- i=391, alt=5, thresh=4.62902e-032, actual=9.04106e-035, err=0
        "1101000101110000001101111100011101", -- i=392, alt=24, thresh=3.15748e-032, actual=6.16695e-035, err=0
        "1101001010000010010000000000110010", -- i=393, alt=4, thresh=2.15162e-032, actual=4.20239e-035, err=5.34553e-051
        "1101001110011111100011110100100010", -- i=394, alt=19, thresh=1.46477e-032, actual=2.86087e-035, err=0
        "1101010011000100011000111110100011", -- i=395, alt=28, thresh=9.96199e-033, actual=1.9457e-035, err=2.67276e-051
        "1101010111001101101011111010010010", -- i=396, alt=3, thresh=6.76861e-033, actual=1.32199e-035, err=2.67276e-051
        "1101011100000100101000000010000010", -- i=397, alt=32, thresh=4.59439e-033, actual=8.97342e-036, err=1.33638e-051
        "1101011111111010010101111100111000", -- i=398, alt=2, thresh=3.11553e-033, actual=6.08503e-036, err=1.33638e-051
        "1101100101000010100111110011100111", -- i=399, alt=13, thresh=2.11063e-033, actual=4.12233e-036, err=0
        "1101101001001010100111111111101111", -- i=400, alt=1, thresh=1.42846e-033, actual=2.78996e-036, err=0
        "1101101101111110000110001111001010", -- i=401, alt=23, thresh=9.65828e-034, actual=1.88638e-036, err=0
        "1101110010011100110100111001011100", -- i=402, alt=18, thresh=6.52389e-034, actual=1.2742e-036, err=0
        "1101110110110110110100100100001011", -- i=403, alt=12, thresh=4.40239e-034, actual=8.59843e-037, err=0
        "1101111011101011000000000011000100", -- i=404, alt=27, thresh=2.96789e-034, actual=5.79665e-037, err=8.35239e-053
        "1101111111101100100111010001111011", -- i=405, alt=31, thresh=1.99885e-034, actual=3.90401e-037, err=0
        "1110000100110100111011011010000000", -- i=406, alt=11, thresh=1.3449e-034, actual=2.62676e-037, err=0
        "1110001000111110101100000000001010", -- i=407, alt=22, thresh=9.04014e-035, actual=1.76565e-037, err=0
        "1110001101111010011101010000001100", -- i=408, alt=17, thresh=6.07066e-035, actual=1.18568e-037, err=0
        "1110010010011101110110101000100011", -- i=409, alt=10, thresh=4.0726e-035, actual=7.9543e-038, err=0
        "1110010110111011011111111011011110", -- i=410, alt=26, thresh=2.7295e-035, actual=5.33106e-038, err=0
        "1110011011110110101001001010010111", -- i=411, alt=30, thresh=1.82756e-035, actual=3.56945e-038, err=5.22024e-054
        "1110011111111000000001100001101110", -- i=412, alt=16, thresh=1.22246e-035, actual=2.38761e-038, err=0
        "1110100101001001000011010110111011", -- i=413, alt=9, thresh=8.16907e-036, actual=1.59552e-038, err=0
        "1110101001100000000111000100111100", -- i=414, alt=21, thresh=5.45364e-036, actual=1.06516e-038, err=1.30506e-054
        "1110101110010101001001100010100111", -- i=415, alt=8, thresh=3.63728e-036, actual=7.10406e-039, err=1.30506e-054
        "1110110011000111010100111101110000", -- i=416, alt=25, thresh=2.42349e-036, actual=4.73339e-039, err=0
        "1110110111011011000100000010000000", -- i=417, alt=15, thresh=1.61318e-036, actual=3.15074e-039, err=6.5253e-055
        "1110111111111111111111111111111111", -- i=418, alt=29, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=419, alt=7, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=420, alt=20, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=421, alt=6, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=422, alt=14, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=423, alt=5, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=424, alt=24, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=425, alt=4, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=426, alt=19, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=427, alt=28, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=428, alt=3, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=429, alt=2, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=430, alt=13, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=431, alt=1, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=432, alt=23, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=433, alt=18, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=434, alt=12, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=435, alt=27, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=436, alt=11, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=437, alt=22, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=438, alt=17, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=439, alt=10, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=440, alt=26, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=441, alt=16, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=442, alt=9, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=443, alt=21, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=444, alt=8, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=445, alt=25, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=446, alt=15, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=447, alt=7, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=448, alt=20, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=449, alt=6, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=450, alt=14, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=451, alt=5, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=452, alt=24, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=453, alt=4, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=454, alt=19, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=455, alt=3, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=456, alt=2, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=457, alt=13, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=458, alt=1, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=459, alt=23, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=460, alt=18, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=461, alt=12, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=462, alt=11, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=463, alt=22, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=464, alt=17, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=465, alt=10, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=466, alt=16, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=467, alt=9, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=468, alt=21, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=469, alt=8, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=470, alt=15, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=471, alt=7, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=472, alt=20, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=473, alt=6, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=474, alt=14, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=475, alt=5, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=476, alt=4, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=477, alt=19, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=478, alt=3, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=479, alt=2, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=480, alt=13, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=481, alt=1, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=482, alt=18, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=483, alt=12, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=484, alt=11, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=485, alt=17, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=486, alt=10, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=487, alt=16, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=488, alt=9, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=489, alt=8, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=490, alt=15, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=491, alt=7, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=492, alt=6, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=493, alt=14, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=494, alt=5, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=495, alt=4, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=496, alt=3, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=497, alt=2, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=498, alt=13, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=499, alt=1, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=500, alt=12, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=501, alt=11, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=502, alt=10, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=503, alt=9, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=504, alt=8, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=505, alt=7, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=506, alt=6, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=507, alt=5, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=508, alt=4, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=509, alt=3, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111", -- i=510, alt=2, thresh=0, actual=0, err=0
        "1110111111111111111111111111111111" -- i=511, alt=1, thresh=0, actual=0, err=0
    );
    attribute rom_style of alias_rom:signal is "block";
    signal c1_alias_thresh_bits : unsigned(67-1 downto 0);
    signal c1_alias_thresh_bits_lo : unsigned(34-1 downto 0);
    signal c1_alias_thresh_bits_lo_d1 : unsigned(34-1 downto 0);
    signal c1_alias_thresh_bits_lo_d2 : unsigned(34-1 downto 0);
    signal c1_alias_thresh_bits_lo_d3 : unsigned(34-1 downto 0);
    signal c1_alias_thresh_bits_hi : unsigned(34-1 downto 0);
    signal c1_alias_thresh_bits_hi_d1 : unsigned(34-1 downto 0);
    signal c1_alias_thresh_bits_hi_d2 : unsigned(34-1 downto 0);
    signal c1_alias_thresh_bits_hi_d3 : unsigned(34-1 downto 0);
    signal c1_alias_index : unsigned(9-1 downto 0);
    signal c1_alias_index_d1 : unsigned(9-1 downto 0);
    signal c1_alias_index_d2 : unsigned(9-1 downto 0);
    signal c1_alias_index_d3 : unsigned(9-1 downto 0);
    signal c2_alias_alt : unsigned(9-1 downto 0);
    signal c2_alias_alt_d1 : unsigned(9-1 downto 0);
    signal c2_alias_index : unsigned(9-1 downto 0);
    signal c2_alias_index_d1 : unsigned(9-1 downto 0);
    signal cltfx_out : std_logic_vector(18-1 downto 0);
    signal cltfx_urng : std_logic_vector(120-1 downto 0);
    signal cltfx_sum_8_1 : signed(15-1 downto 0);
    signal cltfx_sum_8_2 : signed(15-1 downto 0);
    signal cltfx_sum_8_3 : signed(15-1 downto 0);
    signal cltfx_sum_8_4 : signed(15-1 downto 0);
    signal cltfx_sum_8_5 : signed(15-1 downto 0);
    signal cltfx_sum_8_6 : signed(15-1 downto 0);
    signal cltfx_sum_8_7 : signed(15-1 downto 0);
    signal cltfx_sum_8_8 : signed(15-1 downto 0);
    signal cltfx_sum_4_1 : signed(16-1 downto 0);
    signal cltfx_sum_4_2 : signed(16-1 downto 0);
    signal cltfx_sum_4_3 : signed(16-1 downto 0);
    signal cltfx_sum_4_4 : signed(16-1 downto 0);
    signal cltfx_sum_2_1 : signed(17-1 downto 0);
    signal cltfx_sum_2_2 : signed(17-1 downto 0);
    signal cltfx_sum_1_1 : signed(18-1 downto 0);
    --Mixture PDF
    signal mixture_pdf_urng : std_logic_vector(300-1 downto 0);
    signal c0_mixture_sign_flag : std_logic;
    signal c1_mixture_sindex : signed(10-1 downto 0);
    signal mixture_pdf_out : std_logic_vector(26-1 downto 0);
begin
--Render glue
    urng : entity work.urng_w300 generic map(W=>300) port map(clk=>iClk,ce=>iCE,load_en=>iLoadEn,load_data=>iLoadData,rng=>iURNG);
    mixture_pdf_urng<=iURNG;
    oRes<=std_logic_vector(mixture_pdf_out);
--Implementation
    --Bernoulli
    bernoulli_fp_cx_exp_urng <= bernoulli_fp_urng(170-1 downto 51);
    bernoulli_fp_c0_exp_thresh <= unsigned(bernoulli_fp_thresh(58-1 downto 51));
    bernoulli_fp_c0_frac_rand <= unsigned(bernoulli_fp_urng(51-1 downto 0));
    bernoulli_fp_c0_frac_thresh <= unsigned(bernoulli_fp_thresh(51-1 downto 0));
    bernoulli_fp_out <= bernoulli_fp_c1_exp_greater or (bernoulli_fp_c1_exp_equal and bernoulli_fp_c1_frac_greater);

    lmz_branch_1_sig <=  to_unsigned(0,7) when bernoulli_fp_cx_exp_urng(0) = '1' else
             to_unsigned(1,7) when bernoulli_fp_cx_exp_urng(1) = '1' else
             to_unsigned(2,7) when bernoulli_fp_cx_exp_urng(2) = '1' else
             to_unsigned(3,7) when bernoulli_fp_cx_exp_urng(3) = '1' else
             to_unsigned(4,7) when bernoulli_fp_cx_exp_urng(4) = '1' else
             to_unsigned(5,7) when bernoulli_fp_cx_exp_urng(5) = '1' else
             to_unsigned(6,7) when bernoulli_fp_cx_exp_urng(6) = '1' else
             to_unsigned(7,7);
    lmz_branch_hit_1_sig <= bernoulli_fp_cx_exp_urng(7 downto 0) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_2_sig <=  to_unsigned(8,7) when bernoulli_fp_cx_exp_urng(8) = '1' else
             to_unsigned(9,7) when bernoulli_fp_cx_exp_urng(9) = '1' else
             to_unsigned(10,7) when bernoulli_fp_cx_exp_urng(10) = '1' else
             to_unsigned(11,7) when bernoulli_fp_cx_exp_urng(11) = '1' else
             to_unsigned(12,7) when bernoulli_fp_cx_exp_urng(12) = '1' else
             to_unsigned(13,7) when bernoulli_fp_cx_exp_urng(13) = '1' else
             to_unsigned(14,7) when bernoulli_fp_cx_exp_urng(14) = '1' else
             to_unsigned(15,7);
    lmz_branch_hit_2_sig <= bernoulli_fp_cx_exp_urng(15 downto 8) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_3_sig <=  to_unsigned(16,7) when bernoulli_fp_cx_exp_urng(16) = '1' else
             to_unsigned(17,7) when bernoulli_fp_cx_exp_urng(17) = '1' else
             to_unsigned(18,7) when bernoulli_fp_cx_exp_urng(18) = '1' else
             to_unsigned(19,7) when bernoulli_fp_cx_exp_urng(19) = '1' else
             to_unsigned(20,7) when bernoulli_fp_cx_exp_urng(20) = '1' else
             to_unsigned(21,7) when bernoulli_fp_cx_exp_urng(21) = '1' else
             to_unsigned(22,7) when bernoulli_fp_cx_exp_urng(22) = '1' else
             to_unsigned(23,7);
    lmz_branch_hit_3_sig <= bernoulli_fp_cx_exp_urng(23 downto 16) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_4_sig <=  to_unsigned(24,7) when bernoulli_fp_cx_exp_urng(24) = '1' else
             to_unsigned(25,7) when bernoulli_fp_cx_exp_urng(25) = '1' else
             to_unsigned(26,7) when bernoulli_fp_cx_exp_urng(26) = '1' else
             to_unsigned(27,7) when bernoulli_fp_cx_exp_urng(27) = '1' else
             to_unsigned(28,7) when bernoulli_fp_cx_exp_urng(28) = '1' else
             to_unsigned(29,7) when bernoulli_fp_cx_exp_urng(29) = '1' else
             to_unsigned(30,7) when bernoulli_fp_cx_exp_urng(30) = '1' else
             to_unsigned(31,7);
    lmz_branch_hit_4_sig <= bernoulli_fp_cx_exp_urng(31 downto 24) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_5_sig <=  to_unsigned(32,7) when bernoulli_fp_cx_exp_urng(32) = '1' else
             to_unsigned(33,7) when bernoulli_fp_cx_exp_urng(33) = '1' else
             to_unsigned(34,7) when bernoulli_fp_cx_exp_urng(34) = '1' else
             to_unsigned(35,7) when bernoulli_fp_cx_exp_urng(35) = '1' else
             to_unsigned(36,7) when bernoulli_fp_cx_exp_urng(36) = '1' else
             to_unsigned(37,7) when bernoulli_fp_cx_exp_urng(37) = '1' else
             to_unsigned(38,7) when bernoulli_fp_cx_exp_urng(38) = '1' else
             to_unsigned(39,7);
    lmz_branch_hit_5_sig <= bernoulli_fp_cx_exp_urng(39 downto 32) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_6_sig <=  to_unsigned(40,7) when bernoulli_fp_cx_exp_urng(40) = '1' else
             to_unsigned(41,7) when bernoulli_fp_cx_exp_urng(41) = '1' else
             to_unsigned(42,7) when bernoulli_fp_cx_exp_urng(42) = '1' else
             to_unsigned(43,7) when bernoulli_fp_cx_exp_urng(43) = '1' else
             to_unsigned(44,7) when bernoulli_fp_cx_exp_urng(44) = '1' else
             to_unsigned(45,7) when bernoulli_fp_cx_exp_urng(45) = '1' else
             to_unsigned(46,7) when bernoulli_fp_cx_exp_urng(46) = '1' else
             to_unsigned(47,7);
    lmz_branch_hit_6_sig <= bernoulli_fp_cx_exp_urng(47 downto 40) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_7_sig <=  to_unsigned(48,7) when bernoulli_fp_cx_exp_urng(48) = '1' else
             to_unsigned(49,7) when bernoulli_fp_cx_exp_urng(49) = '1' else
             to_unsigned(50,7) when bernoulli_fp_cx_exp_urng(50) = '1' else
             to_unsigned(51,7) when bernoulli_fp_cx_exp_urng(51) = '1' else
             to_unsigned(52,7) when bernoulli_fp_cx_exp_urng(52) = '1' else
             to_unsigned(53,7) when bernoulli_fp_cx_exp_urng(53) = '1' else
             to_unsigned(54,7) when bernoulli_fp_cx_exp_urng(54) = '1' else
             to_unsigned(55,7);
    lmz_branch_hit_7_sig <= bernoulli_fp_cx_exp_urng(55 downto 48) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_8_sig <=  to_unsigned(56,7) when bernoulli_fp_cx_exp_urng(56) = '1' else
             to_unsigned(57,7) when bernoulli_fp_cx_exp_urng(57) = '1' else
             to_unsigned(58,7) when bernoulli_fp_cx_exp_urng(58) = '1' else
             to_unsigned(59,7) when bernoulli_fp_cx_exp_urng(59) = '1' else
             to_unsigned(60,7) when bernoulli_fp_cx_exp_urng(60) = '1' else
             to_unsigned(61,7) when bernoulli_fp_cx_exp_urng(61) = '1' else
             to_unsigned(62,7) when bernoulli_fp_cx_exp_urng(62) = '1' else
             to_unsigned(63,7);
    lmz_branch_hit_8_sig <= bernoulli_fp_cx_exp_urng(63 downto 56) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_9_sig <=  to_unsigned(64,7) when bernoulli_fp_cx_exp_urng(64) = '1' else
             to_unsigned(65,7) when bernoulli_fp_cx_exp_urng(65) = '1' else
             to_unsigned(66,7) when bernoulli_fp_cx_exp_urng(66) = '1' else
             to_unsigned(67,7) when bernoulli_fp_cx_exp_urng(67) = '1' else
             to_unsigned(68,7) when bernoulli_fp_cx_exp_urng(68) = '1' else
             to_unsigned(69,7) when bernoulli_fp_cx_exp_urng(69) = '1' else
             to_unsigned(70,7) when bernoulli_fp_cx_exp_urng(70) = '1' else
             to_unsigned(71,7);
    lmz_branch_hit_9_sig <= bernoulli_fp_cx_exp_urng(71 downto 64) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_10_sig <=  to_unsigned(72,7) when bernoulli_fp_cx_exp_urng(72) = '1' else
             to_unsigned(73,7) when bernoulli_fp_cx_exp_urng(73) = '1' else
             to_unsigned(74,7) when bernoulli_fp_cx_exp_urng(74) = '1' else
             to_unsigned(75,7) when bernoulli_fp_cx_exp_urng(75) = '1' else
             to_unsigned(76,7) when bernoulli_fp_cx_exp_urng(76) = '1' else
             to_unsigned(77,7) when bernoulli_fp_cx_exp_urng(77) = '1' else
             to_unsigned(78,7) when bernoulli_fp_cx_exp_urng(78) = '1' else
             to_unsigned(79,7);
    lmz_branch_hit_10_sig <= bernoulli_fp_cx_exp_urng(79 downto 72) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_11_sig <=  to_unsigned(80,7) when bernoulli_fp_cx_exp_urng(80) = '1' else
             to_unsigned(81,7) when bernoulli_fp_cx_exp_urng(81) = '1' else
             to_unsigned(82,7) when bernoulli_fp_cx_exp_urng(82) = '1' else
             to_unsigned(83,7) when bernoulli_fp_cx_exp_urng(83) = '1' else
             to_unsigned(84,7) when bernoulli_fp_cx_exp_urng(84) = '1' else
             to_unsigned(85,7) when bernoulli_fp_cx_exp_urng(85) = '1' else
             to_unsigned(86,7) when bernoulli_fp_cx_exp_urng(86) = '1' else
             to_unsigned(87,7);
    lmz_branch_hit_11_sig <= bernoulli_fp_cx_exp_urng(87 downto 80) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_12_sig <=  to_unsigned(88,7) when bernoulli_fp_cx_exp_urng(88) = '1' else
             to_unsigned(89,7) when bernoulli_fp_cx_exp_urng(89) = '1' else
             to_unsigned(90,7) when bernoulli_fp_cx_exp_urng(90) = '1' else
             to_unsigned(91,7) when bernoulli_fp_cx_exp_urng(91) = '1' else
             to_unsigned(92,7) when bernoulli_fp_cx_exp_urng(92) = '1' else
             to_unsigned(93,7) when bernoulli_fp_cx_exp_urng(93) = '1' else
             to_unsigned(94,7) when bernoulli_fp_cx_exp_urng(94) = '1' else
             to_unsigned(95,7);
    lmz_branch_hit_12_sig <= bernoulli_fp_cx_exp_urng(95 downto 88) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_13_sig <=  to_unsigned(96,7) when bernoulli_fp_cx_exp_urng(96) = '1' else
             to_unsigned(97,7) when bernoulli_fp_cx_exp_urng(97) = '1' else
             to_unsigned(98,7) when bernoulli_fp_cx_exp_urng(98) = '1' else
             to_unsigned(99,7) when bernoulli_fp_cx_exp_urng(99) = '1' else
             to_unsigned(100,7) when bernoulli_fp_cx_exp_urng(100) = '1' else
             to_unsigned(101,7) when bernoulli_fp_cx_exp_urng(101) = '1' else
             to_unsigned(102,7) when bernoulli_fp_cx_exp_urng(102) = '1' else
             to_unsigned(103,7);
    lmz_branch_hit_13_sig <= bernoulli_fp_cx_exp_urng(103 downto 96) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_14_sig <=  to_unsigned(104,7) when bernoulli_fp_cx_exp_urng(104) = '1' else
             to_unsigned(105,7) when bernoulli_fp_cx_exp_urng(105) = '1' else
             to_unsigned(106,7) when bernoulli_fp_cx_exp_urng(106) = '1' else
             to_unsigned(107,7) when bernoulli_fp_cx_exp_urng(107) = '1' else
             to_unsigned(108,7) when bernoulli_fp_cx_exp_urng(108) = '1' else
             to_unsigned(109,7) when bernoulli_fp_cx_exp_urng(109) = '1' else
             to_unsigned(110,7) when bernoulli_fp_cx_exp_urng(110) = '1' else
             to_unsigned(111,7);
    lmz_branch_hit_14_sig <= bernoulli_fp_cx_exp_urng(111 downto 104) /= std_logic_vector(to_unsigned(0,8));

    lmz_branch_15_sig <=  to_unsigned(112,7) when bernoulli_fp_cx_exp_urng(112) = '1' else
             to_unsigned(113,7) when bernoulli_fp_cx_exp_urng(113) = '1' else
             to_unsigned(114,7) when bernoulli_fp_cx_exp_urng(114) = '1' else
             to_unsigned(115,7) when bernoulli_fp_cx_exp_urng(115) = '1' else
             to_unsigned(116,7) when bernoulli_fp_cx_exp_urng(116) = '1' else
             to_unsigned(117,7) when bernoulli_fp_cx_exp_urng(117) = '1' else
             to_unsigned(118,7);
    lmz_branch_hit_15_sig <= bernoulli_fp_cx_exp_urng(118 downto 112) /= std_logic_vector(to_unsigned(0,7));
    bernoulli_fp_cx_exp_rand <=
        lmz_branch_1 when lmz_branch_hit_1 else
        lmz_branch_2 when lmz_branch_hit_2 else
        lmz_branch_3 when lmz_branch_hit_3 else
        lmz_branch_4 when lmz_branch_hit_4 else
        lmz_branch_5 when lmz_branch_hit_5 else
        lmz_branch_6 when lmz_branch_hit_6 else
        lmz_branch_7 when lmz_branch_hit_7 else
        lmz_branch_8 when lmz_branch_hit_8 else
        lmz_branch_9 when lmz_branch_hit_9 else
        lmz_branch_10 when lmz_branch_hit_10 else
        lmz_branch_11 when lmz_branch_hit_11 else
        lmz_branch_12 when lmz_branch_hit_12 else
        lmz_branch_13 when lmz_branch_hit_13 else
        lmz_branch_14 when lmz_branch_hit_14 else
        lmz_branch_15 when lmz_branch_hit_15 else
        to_unsigned(119,7);

    bernoulli_fp_c0_exp_rand <= bernoulli_fp_c0_exp_rand_d2;
    --Alias table
    c0_alias_index <= unsigned(alias_table_urng(9-1 downto 0));
    bernoulli_fp_urng <= alias_table_urng(179-1 downto 9);
    bernoulli_fp_thresh <= c1_alias_thresh_bits(67-1 downto 9);
    c1_alias_thresh_bits <= c1_alias_thresh_bits_lo&resize(c1_alias_thresh_bits_hi,33);

    c1_alias_thresh_bits_hi <= c1_alias_thresh_bits_hi_d3;

    c1_alias_thresh_bits_lo <= c1_alias_thresh_bits_lo_d3;

    c1_alias_index <= c1_alias_index_d3;

    c2_alias_alt <= c2_alias_alt_d1;

    c2_alias_index <= c2_alias_index_d1;

    cltfx_sum_8_1 <= signed(cltfx_urng(15-1 downto 0));
    cltfx_sum_8_2 <= signed(cltfx_urng(30-1 downto 15));
    cltfx_sum_8_3 <= signed(cltfx_urng(45-1 downto 30));
    cltfx_sum_8_4 <= signed(cltfx_urng(60-1 downto 45));
    cltfx_sum_8_5 <= signed(cltfx_urng(75-1 downto 60));
    cltfx_sum_8_6 <= signed(cltfx_urng(90-1 downto 75));
    cltfx_sum_8_7 <= signed(cltfx_urng(105-1 downto 90));
    cltfx_sum_8_8 <= signed(cltfx_urng(120-1 downto 105));
    cltfx_out<= std_logic_vector(cltfx_sum_1_1);
    --Alias table
    alias_table_urng <= mixture_pdf_urng(179-1 downto 0);
    cltfx_urng <= mixture_pdf_urng(299-1 downto 179);
    c0_mixture_sign_flag <= mixture_pdf_urng(299);
process(iClk) begin if(rising_edge(iClk)) then if(iCE='1') then
    --Bernoulli

    lmz_branch_1 <= lmz_branch_1_sig;
    lmz_branch_hit_1 <= lmz_branch_hit_1_sig;
    lmz_branch_2 <= lmz_branch_2_sig;
    lmz_branch_hit_2 <= lmz_branch_hit_2_sig;
    lmz_branch_3 <= lmz_branch_3_sig;
    lmz_branch_hit_3 <= lmz_branch_hit_3_sig;
    lmz_branch_4 <= lmz_branch_4_sig;
    lmz_branch_hit_4 <= lmz_branch_hit_4_sig;
    lmz_branch_5 <= lmz_branch_5_sig;
    lmz_branch_hit_5 <= lmz_branch_hit_5_sig;
    lmz_branch_6 <= lmz_branch_6_sig;
    lmz_branch_hit_6 <= lmz_branch_hit_6_sig;
    lmz_branch_7 <= lmz_branch_7_sig;
    lmz_branch_hit_7 <= lmz_branch_hit_7_sig;
    lmz_branch_8 <= lmz_branch_8_sig;
    lmz_branch_hit_8 <= lmz_branch_hit_8_sig;
    lmz_branch_9 <= lmz_branch_9_sig;
    lmz_branch_hit_9 <= lmz_branch_hit_9_sig;
    lmz_branch_10 <= lmz_branch_10_sig;
    lmz_branch_hit_10 <= lmz_branch_hit_10_sig;
    lmz_branch_11 <= lmz_branch_11_sig;
    lmz_branch_hit_11 <= lmz_branch_hit_11_sig;
    lmz_branch_12 <= lmz_branch_12_sig;
    lmz_branch_hit_12 <= lmz_branch_hit_12_sig;
    lmz_branch_13 <= lmz_branch_13_sig;
    lmz_branch_hit_13 <= lmz_branch_hit_13_sig;
    lmz_branch_14 <= lmz_branch_14_sig;
    lmz_branch_hit_14 <= lmz_branch_hit_14_sig;
    lmz_branch_15 <= lmz_branch_15_sig;
    lmz_branch_hit_15 <= lmz_branch_hit_15_sig;

    bernoulli_fp_c0_exp_rand_d1 <= bernoulli_fp_cx_exp_rand;
    bernoulli_fp_c0_exp_rand_d2 <= bernoulli_fp_c0_exp_rand_d1;
    bernoulli_fp_c1_exp_greater <= bernoulli_fp_c0_exp_rand > bernoulli_fp_c0_exp_thresh;
    bernoulli_fp_c1_exp_equal <= bernoulli_fp_c0_exp_rand = bernoulli_fp_c0_exp_thresh;
    bernoulli_fp_c1_frac_greater <= bernoulli_fp_c0_frac_rand > bernoulli_fp_c0_frac_thresh;
    --Alias table

    c1_alias_thresh_bits_hi_d1 <= alias_rom(to_integer('0'&c0_alias_index));
    c1_alias_thresh_bits_hi_d2 <= c1_alias_thresh_bits_hi_d1;
    c1_alias_thresh_bits_hi_d3 <= c1_alias_thresh_bits_hi_d2;

    c1_alias_thresh_bits_lo_d1 <= alias_rom(to_integer('1'&c0_alias_index));
    c1_alias_thresh_bits_lo_d2 <= c1_alias_thresh_bits_lo_d1;
    c1_alias_thresh_bits_lo_d3 <= c1_alias_thresh_bits_lo_d2;

    c1_alias_index_d1 <= c0_alias_index;
    c1_alias_index_d2 <= c1_alias_index_d1;
    c1_alias_index_d3 <= c1_alias_index_d2;

    c2_alias_alt_d1 <= c1_alias_thresh_bits(9-1 downto 0);

    c2_alias_index_d1 <= c1_alias_index;
    if bernoulli_fp_out then
        alias_table_out <= c2_alias_index;
    else
        alias_table_out <= c2_alias_alt;
    end if;

    cltfx_sum_4_1 <= resize(cltfx_sum_8_2,16) - resize(cltfx_sum_8_1,16);
    cltfx_sum_4_2 <= resize(cltfx_sum_8_4,16) - resize(cltfx_sum_8_3,16);
    cltfx_sum_4_3 <= resize(cltfx_sum_8_6,16) - resize(cltfx_sum_8_5,16);
    cltfx_sum_4_4 <= resize(cltfx_sum_8_8,16) - resize(cltfx_sum_8_7,16);
    cltfx_sum_2_1 <= resize(cltfx_sum_4_2,17) - resize(cltfx_sum_4_1,17);
    cltfx_sum_2_2 <= resize(cltfx_sum_4_4,17) - resize(cltfx_sum_4_3,17);
    cltfx_sum_1_1 <= resize(cltfx_sum_2_2,18) - resize(cltfx_sum_2_1,18);
    --Alias table
    if c0_mixture_sign_flag='1' then
        c1_mixture_sindex <= signed(resize(unsigned(alias_table_out),10));
    else
        c1_mixture_sindex <= -signed(resize(unsigned(alias_table_out),10));
    end if;
    mixture_pdf_out <= std_logic_vector(resize(signed(cltfx_out),26) + ((resize(c1_mixture_sindex,26) sll 15)));
end if; end if; end process;
end RTL;
