
library ieee;
use ieee.std_logic_1164.all;

entity rng_n234_r234_t5_k0_s3206 is
  port(
    clk:in std_logic;
    ce:in std_logic;
    mode:in std_logic;
    s_in:in std_logic;
    s_out:out std_logic;
    rng:out std_logic_vector(233 downto 0)
  );
end rng_n234_r234_t5_k0_s3206;

architecture RTL of rng_n234_r234_t5_k0_s3206 is
  signal fifo_out, r_out:std_logic_vector(233 downto 0) := (others=>'1');
begin
  rng(0) <= r_out(232);
  rng(1) <= r_out(22);
  rng(2) <= r_out(207);
  rng(3) <= r_out(11);
  rng(4) <= r_out(3);
  rng(5) <= r_out(14);
  rng(6) <= r_out(191);
  rng(7) <= r_out(156);
  rng(8) <= r_out(117);
  rng(9) <= r_out(37);
  rng(10) <= r_out(38);
  rng(11) <= r_out(40);
  rng(12) <= r_out(44);
  rng(13) <= r_out(119);
  rng(14) <= r_out(66);
  rng(15) <= r_out(181);
  rng(16) <= r_out(176);
  rng(17) <= r_out(65);
  rng(18) <= r_out(5);
  rng(19) <= r_out(233);
  rng(20) <= r_out(16);
  rng(21) <= r_out(141);
  rng(22) <= r_out(1);
  rng(23) <= r_out(32);
  rng(24) <= r_out(228);
  rng(25) <= r_out(157);
  rng(26) <= r_out(70);
  rng(27) <= r_out(53);
  rng(28) <= r_out(116);
  rng(29) <= r_out(204);
  rng(30) <= r_out(85);
  rng(31) <= r_out(35);
  rng(32) <= r_out(159);
  rng(33) <= r_out(106);
  rng(34) <= r_out(222);
  rng(35) <= r_out(166);
  rng(36) <= r_out(122);
  rng(37) <= r_out(86);
  rng(38) <= r_out(81);
  rng(39) <= r_out(50);
  rng(40) <= r_out(225);
  rng(41) <= r_out(9);
  rng(42) <= r_out(109);
  rng(43) <= r_out(138);
  rng(44) <= r_out(77);
  rng(45) <= r_out(148);
  rng(46) <= r_out(91);
  rng(47) <= r_out(76);
  rng(48) <= r_out(127);
  rng(49) <= r_out(188);
  rng(50) <= r_out(60);
  rng(51) <= r_out(190);
  rng(52) <= r_out(193);
  rng(53) <= r_out(113);
  rng(54) <= r_out(226);
  rng(55) <= r_out(97);
  rng(56) <= r_out(154);
  rng(57) <= r_out(72);
  rng(58) <= r_out(47);
  rng(59) <= r_out(203);
  rng(60) <= r_out(135);
  rng(61) <= r_out(223);
  rng(62) <= r_out(105);
  rng(63) <= r_out(183);
  rng(64) <= r_out(147);
  rng(65) <= r_out(15);
  rng(66) <= r_out(199);
  rng(67) <= r_out(187);
  rng(68) <= r_out(87);
  rng(69) <= r_out(96);
  rng(70) <= r_out(214);
  rng(71) <= r_out(94);
  rng(72) <= r_out(175);
  rng(73) <= r_out(151);
  rng(74) <= r_out(230);
  rng(75) <= r_out(196);
  rng(76) <= r_out(150);
  rng(77) <= r_out(205);
  rng(78) <= r_out(123);
  rng(79) <= r_out(200);
  rng(80) <= r_out(144);
  rng(81) <= r_out(213);
  rng(82) <= r_out(90);
  rng(83) <= r_out(59);
  rng(84) <= r_out(18);
  rng(85) <= r_out(163);
  rng(86) <= r_out(218);
  rng(87) <= r_out(126);
  rng(88) <= r_out(224);
  rng(89) <= r_out(45);
  rng(90) <= r_out(110);
  rng(91) <= r_out(78);
  rng(92) <= r_out(24);
  rng(93) <= r_out(136);
  rng(94) <= r_out(12);
  rng(95) <= r_out(92);
  rng(96) <= r_out(67);
  rng(97) <= r_out(71);
  rng(98) <= r_out(186);
  rng(99) <= r_out(129);
  rng(100) <= r_out(130);
  rng(101) <= r_out(104);
  rng(102) <= r_out(145);
  rng(103) <= r_out(4);
  rng(104) <= r_out(158);
  rng(105) <= r_out(137);
  rng(106) <= r_out(101);
  rng(107) <= r_out(20);
  rng(108) <= r_out(68);
  rng(109) <= r_out(114);
  rng(110) <= r_out(133);
  rng(111) <= r_out(179);
  rng(112) <= r_out(197);
  rng(113) <= r_out(167);
  rng(114) <= r_out(206);
  rng(115) <= r_out(182);
  rng(116) <= r_out(189);
  rng(117) <= r_out(17);
  rng(118) <= r_out(131);
  rng(119) <= r_out(140);
  rng(120) <= r_out(146);
  rng(121) <= r_out(30);
  rng(122) <= r_out(69);
  rng(123) <= r_out(62);
  rng(124) <= r_out(100);
  rng(125) <= r_out(10);
  rng(126) <= r_out(171);
  rng(127) <= r_out(219);
  rng(128) <= r_out(209);
  rng(129) <= r_out(52);
  rng(130) <= r_out(98);
  rng(131) <= r_out(46);
  rng(132) <= r_out(210);
  rng(133) <= r_out(192);
  rng(134) <= r_out(198);
  rng(135) <= r_out(64);
  rng(136) <= r_out(115);
  rng(137) <= r_out(211);
  rng(138) <= r_out(95);
  rng(139) <= r_out(83);
  rng(140) <= r_out(33);
  rng(141) <= r_out(194);
  rng(142) <= r_out(93);
  rng(143) <= r_out(103);
  rng(144) <= r_out(42);
  rng(145) <= r_out(220);
  rng(146) <= r_out(27);
  rng(147) <= r_out(23);
  rng(148) <= r_out(217);
  rng(149) <= r_out(143);
  rng(150) <= r_out(177);
  rng(151) <= r_out(112);
  rng(152) <= r_out(216);
  rng(153) <= r_out(229);
  rng(154) <= r_out(162);
  rng(155) <= r_out(184);
  rng(156) <= r_out(155);
  rng(157) <= r_out(202);
  rng(158) <= r_out(124);
  rng(159) <= r_out(99);
  rng(160) <= r_out(13);
  rng(161) <= r_out(55);
  rng(162) <= r_out(26);
  rng(163) <= r_out(142);
  rng(164) <= r_out(29);
  rng(165) <= r_out(132);
  rng(166) <= r_out(121);
  rng(167) <= r_out(84);
  rng(168) <= r_out(153);
  rng(169) <= r_out(172);
  rng(170) <= r_out(80);
  rng(171) <= r_out(231);
  rng(172) <= r_out(134);
  rng(173) <= r_out(41);
  rng(174) <= r_out(128);
  rng(175) <= r_out(170);
  rng(176) <= r_out(21);
  rng(177) <= r_out(102);
  rng(178) <= r_out(208);
  rng(179) <= r_out(185);
  rng(180) <= r_out(43);
  rng(181) <= r_out(178);
  rng(182) <= r_out(168);
  rng(183) <= r_out(25);
  rng(184) <= r_out(49);
  rng(185) <= r_out(221);
  rng(186) <= r_out(8);
  rng(187) <= r_out(139);
  rng(188) <= r_out(73);
  rng(189) <= r_out(79);
  rng(190) <= r_out(120);
  rng(191) <= r_out(58);
  rng(192) <= r_out(108);
  rng(193) <= r_out(180);
  rng(194) <= r_out(82);
  rng(195) <= r_out(164);
  rng(196) <= r_out(39);
  rng(197) <= r_out(215);
  rng(198) <= r_out(111);
  rng(199) <= r_out(0);
  rng(200) <= r_out(149);
  rng(201) <= r_out(28);
  rng(202) <= r_out(2);
  rng(203) <= r_out(89);
  rng(204) <= r_out(227);
  rng(205) <= r_out(201);
  rng(206) <= r_out(118);
  rng(207) <= r_out(195);
  rng(208) <= r_out(169);
  rng(209) <= r_out(161);
  rng(210) <= r_out(174);
  rng(211) <= r_out(36);
  rng(212) <= r_out(75);
  rng(213) <= r_out(7);
  rng(214) <= r_out(107);
  rng(215) <= r_out(6);
  rng(216) <= r_out(48);
  rng(217) <= r_out(61);
  rng(218) <= r_out(54);
  rng(219) <= r_out(56);
  rng(220) <= r_out(19);
  rng(221) <= r_out(63);
  rng(222) <= r_out(88);
  rng(223) <= r_out(51);
  rng(224) <= r_out(173);
  rng(225) <= r_out(34);
  rng(226) <= r_out(31);
  rng(227) <= r_out(74);
  rng(228) <= r_out(125);
  rng(229) <= r_out(165);
  rng(230) <= r_out(152);
  rng(231) <= r_out(212);
  rng(232) <= r_out(57);
  rng(233) <= r_out(160);
  s_out <= fifo_out(28);
  regs : process(clk) begin
    if(rising_edge(clk)) then if(ce='1') then
      r_out(0)<=(mode and fifo_out(0)) or ((not mode) and ('0' xor fifo_out(0) xor fifo_out(18) xor fifo_out(32) xor fifo_out(40) xor fifo_out(219)));
      r_out(1)<=(mode and fifo_out(1)) or ((not mode) and ('0' xor fifo_out(1) xor fifo_out(111) xor fifo_out(157) xor fifo_out(174) xor fifo_out(185)));
      r_out(2)<=(mode and fifo_out(2)) or ((not mode) and ('0' xor fifo_out(2) xor fifo_out(80) xor fifo_out(134) xor fifo_out(171) xor fifo_out(190)));
      r_out(3)<=(mode and fifo_out(3)) or ((not mode) and ('0' xor fifo_out(3) xor fifo_out(24) xor fifo_out(36) xor fifo_out(49) xor fifo_out(58)));
      r_out(4)<=(mode and fifo_out(4)) or ((not mode) and ('0' xor fifo_out(4) xor fifo_out(39) xor fifo_out(83) xor fifo_out(130) xor fifo_out(220)));
      r_out(5)<=(mode and fifo_out(5)) or ((not mode) and ('0' xor fifo_out(5) xor fifo_out(43) xor fifo_out(62) xor fifo_out(147) xor fifo_out(200)));
      r_out(6)<=(mode and fifo_out(6)) or ((not mode) and ('0' xor fifo_out(6) xor fifo_out(116) xor fifo_out(121) xor fifo_out(209) xor fifo_out(228)));
      r_out(7)<=(mode and fifo_out(7)) or ((not mode) and ('0' xor fifo_out(7) xor fifo_out(50) xor fifo_out(137) xor fifo_out(213) xor fifo_out(226)));
      r_out(8)<=(mode and fifo_out(8)) or ((not mode) and ('0' xor fifo_out(3) xor fifo_out(8) xor fifo_out(176) xor fifo_out(196) xor fifo_out(210)));
      r_out(9)<=(mode and fifo_out(9)) or ((not mode) and ('0' xor fifo_out(9) xor fifo_out(28) xor fifo_out(62) xor fifo_out(86) xor fifo_out(207)));
      r_out(10)<=(mode and fifo_out(10)) or ((not mode) and ('0' xor fifo_out(10) xor fifo_out(55) xor fifo_out(61) xor fifo_out(97) xor fifo_out(152)));
      r_out(11)<=(mode and fifo_out(11)) or ((not mode) and ('0' xor fifo_out(11) xor fifo_out(23) xor fifo_out(77) xor fifo_out(175) xor fifo_out(232)));
      r_out(12)<=(mode and fifo_out(12)) or ((not mode) and ('0' xor fifo_out(12) xor fifo_out(88) xor fifo_out(108) xor fifo_out(141) xor fifo_out(184)));
      r_out(13)<=(mode and fifo_out(13)) or ((not mode) and ('0' xor fifo_out(13) xor fifo_out(99) xor fifo_out(154) xor fifo_out(171) xor fifo_out(185)));
      r_out(14)<=(mode and fifo_out(14)) or ((not mode) and ('0' xor fifo_out(14) xor fifo_out(15) xor fifo_out(129) xor fifo_out(219) xor fifo_out(232)));
      r_out(15)<=(mode and fifo_out(15)) or ((not mode) and ('0' xor fifo_out(15) xor fifo_out(41) xor fifo_out(146) xor fifo_out(152) xor fifo_out(218)));
      r_out(16)<=(mode and fifo_out(16)) or ((not mode) and ('0' xor fifo_out(16) xor fifo_out(50) xor fifo_out(58) xor fifo_out(192) xor fifo_out(199)));
      r_out(17)<=(mode and fifo_out(17)) or ((not mode) and ('0' xor fifo_out(17) xor fifo_out(54) xor fifo_out(108) xor fifo_out(153) xor fifo_out(206)));
      r_out(18)<=(mode and fifo_out(18)) or ((not mode) and ('0' xor fifo_out(9) xor fifo_out(18) xor fifo_out(130) xor fifo_out(198) xor fifo_out(225)));
      r_out(19)<=(mode and fifo_out(19)) or ((not mode) and ('0' xor fifo_out(19) xor fifo_out(69) xor fifo_out(83) xor fifo_out(122) xor fifo_out(178)));
      r_out(20)<=(mode and fifo_out(20)) or ((not mode) and ('0' xor fifo_out(20) xor fifo_out(48) xor fifo_out(80) xor fifo_out(200) xor fifo_out(214)));
      r_out(21)<=(mode and fifo_out(21)) or ((not mode) and ('0' xor fifo_out(21) xor fifo_out(29) xor fifo_out(146) xor fifo_out(194)));
      r_out(22)<=(mode and fifo_out(22)) or ((not mode) and ('0' xor fifo_out(6) xor fifo_out(22) xor fifo_out(74) xor fifo_out(89) xor fifo_out(166)));
      r_out(23)<=(mode and fifo_out(23)) or ((not mode) and ('0' xor fifo_out(23) xor fifo_out(33) xor fifo_out(35) xor fifo_out(191) xor fifo_out(209)));
      r_out(24)<=(mode and fifo_out(24)) or ((not mode) and ('0' xor fifo_out(3) xor fifo_out(24) xor fifo_out(45) xor fifo_out(76) xor fifo_out(161)));
      r_out(25)<=(mode and fifo_out(25)) or ((not mode) and ('0' xor fifo_out(25) xor fifo_out(38) xor fifo_out(60) xor fifo_out(165) xor fifo_out(206)));
      r_out(26)<=(mode and fifo_out(26)) or ((not mode) and ('0' xor fifo_out(26) xor fifo_out(54) xor fifo_out(117) xor fifo_out(155) xor fifo_out(202)));
      r_out(27)<=(mode and fifo_out(27)) or ((not mode) and ('0' xor fifo_out(1) xor fifo_out(21) xor fifo_out(27) xor fifo_out(64) xor fifo_out(164)));
      r_out(28)<=(mode and s_in) or ((not mode) and ('0' xor fifo_out(28) xor fifo_out(52) xor fifo_out(84) xor fifo_out(132)));
      r_out(29)<=(mode and fifo_out(29)) or ((not mode) and ('0' xor fifo_out(29) xor fifo_out(65) xor fifo_out(88) xor fifo_out(131) xor fifo_out(158)));
      r_out(30)<=(mode and fifo_out(30)) or ((not mode) and ('0' xor fifo_out(30) xor fifo_out(143) xor fifo_out(192) xor fifo_out(225) xor fifo_out(226)));
      r_out(31)<=(mode and fifo_out(31)) or ((not mode) and ('0' xor fifo_out(31) xor fifo_out(46) xor fifo_out(59) xor fifo_out(112) xor fifo_out(122)));
      r_out(32)<=(mode and fifo_out(32)) or ((not mode) and ('0' xor fifo_out(17) xor fifo_out(32) xor fifo_out(58) xor fifo_out(136) xor fifo_out(189)));
      r_out(33)<=(mode and fifo_out(33)) or ((not mode) and ('0' xor fifo_out(33) xor fifo_out(128) xor fifo_out(186) xor fifo_out(201) xor fifo_out(215)));
      r_out(34)<=(mode and fifo_out(34)) or ((not mode) and ('0' xor fifo_out(34) xor fifo_out(146) xor fifo_out(149) xor fifo_out(184) xor fifo_out(186)));
      r_out(35)<=(mode and fifo_out(35)) or ((not mode) and ('0' xor fifo_out(21) xor fifo_out(31) xor fifo_out(35) xor fifo_out(194) xor fifo_out(216)));
      r_out(36)<=(mode and fifo_out(36)) or ((not mode) and ('0' xor fifo_out(13) xor fifo_out(17) xor fifo_out(22) xor fifo_out(36) xor fifo_out(109)));
      r_out(37)<=(mode and fifo_out(37)) or ((not mode) and ('0' xor fifo_out(9) xor fifo_out(37) xor fifo_out(82) xor fifo_out(148) xor fifo_out(177)));
      r_out(38)<=(mode and fifo_out(38)) or ((not mode) and ('0' xor fifo_out(12) xor fifo_out(38) xor fifo_out(51) xor fifo_out(66) xor fifo_out(213)));
      r_out(39)<=(mode and fifo_out(39)) or ((not mode) and ('0' xor fifo_out(233) xor fifo_out(39) xor fifo_out(57) xor fifo_out(79) xor fifo_out(152)));
      r_out(40)<=(mode and fifo_out(40)) or ((not mode) and ('0' xor fifo_out(27) xor fifo_out(33) xor fifo_out(40) xor fifo_out(75) xor fifo_out(134)));
      r_out(41)<=(mode and fifo_out(41)) or ((not mode) and ('0' xor fifo_out(41) xor fifo_out(47) xor fifo_out(74) xor fifo_out(93) xor fifo_out(208)));
      r_out(42)<=(mode and fifo_out(42)) or ((not mode) and ('0' xor fifo_out(42) xor fifo_out(103) xor fifo_out(113) xor fifo_out(203) xor fifo_out(207)));
      r_out(43)<=(mode and fifo_out(43)) or ((not mode) and ('0' xor fifo_out(7) xor fifo_out(13) xor fifo_out(43) xor fifo_out(102) xor fifo_out(158)));
      r_out(44)<=(mode and fifo_out(44)) or ((not mode) and ('0' xor fifo_out(44) xor fifo_out(59) xor fifo_out(85) xor fifo_out(129) xor fifo_out(206)));
      r_out(45)<=(mode and fifo_out(45)) or ((not mode) and ('0' xor fifo_out(27) xor fifo_out(45) xor fifo_out(229) xor fifo_out(231) xor fifo_out(232)));
      r_out(46)<=(mode and fifo_out(46)) or ((not mode) and ('0' xor fifo_out(9) xor fifo_out(46) xor fifo_out(131) xor fifo_out(141) xor fifo_out(197)));
      r_out(47)<=(mode and fifo_out(47)) or ((not mode) and ('0' xor fifo_out(17) xor fifo_out(42) xor fifo_out(47) xor fifo_out(77) xor fifo_out(85)));
      r_out(48)<=(mode and fifo_out(48)) or ((not mode) and ('0' xor fifo_out(48) xor fifo_out(110) xor fifo_out(164) xor fifo_out(221) xor fifo_out(225)));
      r_out(49)<=(mode and fifo_out(49)) or ((not mode) and ('0' xor fifo_out(49) xor fifo_out(86) xor fifo_out(94) xor fifo_out(123) xor fifo_out(218)));
      r_out(50)<=(mode and fifo_out(50)) or ((not mode) and ('0' xor fifo_out(50) xor fifo_out(52) xor fifo_out(73) xor fifo_out(226) xor fifo_out(227)));
      r_out(51)<=(mode and fifo_out(51)) or ((not mode) and ('0' xor fifo_out(23) xor fifo_out(51) xor fifo_out(67) xor fifo_out(84) xor fifo_out(199)));
      r_out(52)<=(mode and fifo_out(52)) or ((not mode) and ('0' xor fifo_out(35) xor fifo_out(52) xor fifo_out(96) xor fifo_out(97) xor fifo_out(124)));
      r_out(53)<=(mode and fifo_out(53)) or ((not mode) and ('0' xor fifo_out(10) xor fifo_out(53) xor fifo_out(54) xor fifo_out(189)));
      r_out(54)<=(mode and fifo_out(54)) or ((not mode) and ('0' xor fifo_out(54) xor fifo_out(111) xor fifo_out(115) xor fifo_out(211) xor fifo_out(217)));
      r_out(55)<=(mode and fifo_out(55)) or ((not mode) and ('0' xor fifo_out(3) xor fifo_out(55) xor fifo_out(68) xor fifo_out(159) xor fifo_out(217)));
      r_out(56)<=(mode and fifo_out(56)) or ((not mode) and ('0' xor fifo_out(6) xor fifo_out(25) xor fifo_out(56) xor fifo_out(222) xor fifo_out(227)));
      r_out(57)<=(mode and fifo_out(57)) or ((not mode) and ('0' xor fifo_out(57) xor fifo_out(105) xor fifo_out(180) xor fifo_out(185) xor fifo_out(207)));
      r_out(58)<=(mode and fifo_out(58)) or ((not mode) and ('0' xor fifo_out(36) xor fifo_out(38) xor fifo_out(56) xor fifo_out(58) xor fifo_out(116)));
      r_out(59)<=(mode and fifo_out(59)) or ((not mode) and ('0' xor fifo_out(59) xor fifo_out(106) xor fifo_out(128) xor fifo_out(167) xor fifo_out(172)));
      r_out(60)<=(mode and fifo_out(60)) or ((not mode) and ('0' xor fifo_out(15) xor fifo_out(26) xor fifo_out(60) xor fifo_out(99) xor fifo_out(221)));
      r_out(61)<=(mode and fifo_out(61)) or ((not mode) and ('0' xor fifo_out(3) xor fifo_out(22) xor fifo_out(61) xor fifo_out(168) xor fifo_out(212)));
      r_out(62)<=(mode and fifo_out(62)) or ((not mode) and ('0' xor fifo_out(40) xor fifo_out(62) xor fifo_out(80) xor fifo_out(182) xor fifo_out(230)));
      r_out(63)<=(mode and fifo_out(63)) or ((not mode) and ('0' xor fifo_out(22) xor fifo_out(38) xor fifo_out(63) xor fifo_out(142) xor fifo_out(199)));
      r_out(64)<=(mode and fifo_out(64)) or ((not mode) and ('0' xor fifo_out(11) xor fifo_out(64) xor fifo_out(79) xor fifo_out(132) xor fifo_out(155)));
      r_out(65)<=(mode and fifo_out(65)) or ((not mode) and ('0' xor fifo_out(13) xor fifo_out(16) xor fifo_out(65) xor fifo_out(144) xor fifo_out(188)));
      r_out(66)<=(mode and fifo_out(66)) or ((not mode) and ('0' xor fifo_out(66) xor fifo_out(136) xor fifo_out(164) xor fifo_out(183) xor fifo_out(188)));
      r_out(67)<=(mode and fifo_out(67)) or ((not mode) and ('0' xor fifo_out(6) xor fifo_out(11) xor fifo_out(67) xor fifo_out(72) xor fifo_out(93)));
      r_out(68)<=(mode and fifo_out(68)) or ((not mode) and ('0' xor fifo_out(68) xor fifo_out(126) xor fifo_out(191) xor fifo_out(222) xor fifo_out(223)));
      r_out(69)<=(mode and fifo_out(69)) or ((not mode) and ('0' xor fifo_out(32) xor fifo_out(58) xor fifo_out(69) xor fifo_out(120) xor fifo_out(139)));
      r_out(70)<=(mode and fifo_out(70)) or ((not mode) and ('0' xor fifo_out(4) xor fifo_out(32) xor fifo_out(48) xor fifo_out(70) xor fifo_out(128)));
      r_out(71)<=(mode and fifo_out(71)) or ((not mode) and ('0' xor fifo_out(15) xor fifo_out(71) xor fifo_out(81) xor fifo_out(205) xor fifo_out(221)));
      r_out(72)<=(mode and fifo_out(72)) or ((not mode) and ('0' xor fifo_out(9) xor fifo_out(24) xor fifo_out(72) xor fifo_out(146) xor fifo_out(218)));
      r_out(73)<=(mode and fifo_out(73)) or ((not mode) and ('0' xor fifo_out(39) xor fifo_out(60) xor fifo_out(64) xor fifo_out(73) xor fifo_out(211)));
      r_out(74)<=(mode and fifo_out(74)) or ((not mode) and ('0' xor fifo_out(61) xor fifo_out(74) xor fifo_out(78) xor fifo_out(126) xor fifo_out(211)));
      r_out(75)<=(mode and fifo_out(75)) or ((not mode) and ('0' xor fifo_out(51) xor fifo_out(75) xor fifo_out(81) xor fifo_out(141) xor fifo_out(153)));
      r_out(76)<=(mode and fifo_out(76)) or ((not mode) and ('0' xor fifo_out(71) xor fifo_out(76) xor fifo_out(91) xor fifo_out(138) xor fifo_out(203)));
      r_out(77)<=(mode and fifo_out(77)) or ((not mode) and ('0' xor fifo_out(11) xor fifo_out(74) xor fifo_out(77) xor fifo_out(196)));
      r_out(78)<=(mode and fifo_out(78)) or ((not mode) and ('0' xor fifo_out(23) xor fifo_out(78) xor fifo_out(130) xor fifo_out(155) xor fifo_out(220)));
      r_out(79)<=(mode and fifo_out(79)) or ((not mode) and ('0' xor fifo_out(5) xor fifo_out(62) xor fifo_out(79) xor fifo_out(130) xor fifo_out(224)));
      r_out(80)<=(mode and fifo_out(80)) or ((not mode) and ('0' xor fifo_out(80) xor fifo_out(97) xor fifo_out(116) xor fifo_out(156) xor fifo_out(204)));
      r_out(81)<=(mode and fifo_out(81)) or ((not mode) and ('0' xor fifo_out(44) xor fifo_out(81) xor fifo_out(113) xor fifo_out(123) xor fifo_out(181)));
      r_out(82)<=(mode and fifo_out(82)) or ((not mode) and ('0' xor fifo_out(25) xor fifo_out(78) xor fifo_out(82) xor fifo_out(99) xor fifo_out(151)));
      r_out(83)<=(mode and fifo_out(83)) or ((not mode) and ('0' xor fifo_out(57) xor fifo_out(70) xor fifo_out(83) xor fifo_out(102) xor fifo_out(212)));
      r_out(84)<=(mode and fifo_out(84)) or ((not mode) and ('0' xor fifo_out(39) xor fifo_out(84) xor fifo_out(132) xor fifo_out(183) xor fifo_out(201)));
      r_out(85)<=(mode and fifo_out(85)) or ((not mode) and ('0' xor fifo_out(34) xor fifo_out(50) xor fifo_out(85) xor fifo_out(121) xor fifo_out(219)));
      r_out(86)<=(mode and fifo_out(86)) or ((not mode) and ('0' xor fifo_out(71) xor fifo_out(86) xor fifo_out(90) xor fifo_out(167) xor fifo_out(192)));
      r_out(87)<=(mode and fifo_out(87)) or ((not mode) and ('0' xor fifo_out(87) xor fifo_out(153) xor fifo_out(154) xor fifo_out(193) xor fifo_out(204)));
      r_out(88)<=(mode and fifo_out(88)) or ((not mode) and ('0' xor fifo_out(31) xor fifo_out(88) xor fifo_out(145) xor fifo_out(202) xor fifo_out(226)));
      r_out(89)<=(mode and fifo_out(89)) or ((not mode) and ('0' xor fifo_out(89) xor fifo_out(101) xor fifo_out(107) xor fifo_out(173) xor fifo_out(189)));
      r_out(90)<=(mode and fifo_out(90)) or ((not mode) and ('0' xor fifo_out(26) xor fifo_out(70) xor fifo_out(90) xor fifo_out(176) xor fifo_out(210)));
      r_out(91)<=(mode and fifo_out(91)) or ((not mode) and ('0' xor fifo_out(16) xor fifo_out(57) xor fifo_out(91) xor fifo_out(108) xor fifo_out(215)));
      r_out(92)<=(mode and fifo_out(92)) or ((not mode) and ('0' xor fifo_out(92) xor fifo_out(116) xor fifo_out(150) xor fifo_out(171) xor fifo_out(205)));
      r_out(93)<=(mode and fifo_out(93)) or ((not mode) and ('0' xor fifo_out(82) xor fifo_out(93) xor fifo_out(96) xor fifo_out(160) xor fifo_out(197)));
      r_out(94)<=(mode and fifo_out(94)) or ((not mode) and ('0' xor fifo_out(94) xor fifo_out(138) xor fifo_out(145) xor fifo_out(169)));
      r_out(95)<=(mode and fifo_out(95)) or ((not mode) and ('0' xor fifo_out(95) xor fifo_out(113) xor fifo_out(154) xor fifo_out(162) xor fifo_out(169)));
      r_out(96)<=(mode and fifo_out(96)) or ((not mode) and ('0' xor fifo_out(30) xor fifo_out(84) xor fifo_out(96) xor fifo_out(140) xor fifo_out(166)));
      r_out(97)<=(mode and fifo_out(97)) or ((not mode) and ('0' xor fifo_out(67) xor fifo_out(97) xor fifo_out(133) xor fifo_out(148) xor fifo_out(194)));
      r_out(98)<=(mode and fifo_out(98)) or ((not mode) and ('0' xor fifo_out(98) xor fifo_out(110) xor fifo_out(120) xor fifo_out(124) xor fifo_out(157)));
      r_out(99)<=(mode and fifo_out(99)) or ((not mode) and ('0' xor fifo_out(8) xor fifo_out(83) xor fifo_out(99) xor fifo_out(169) xor fifo_out(191)));
      r_out(100)<=(mode and fifo_out(100)) or ((not mode) and ('0' xor fifo_out(34) xor fifo_out(81) xor fifo_out(100) xor fifo_out(137) xor fifo_out(208)));
      r_out(101)<=(mode and fifo_out(101)) or ((not mode) and ('0' xor fifo_out(47) xor fifo_out(101) xor fifo_out(126) xor fifo_out(165) xor fifo_out(198)));
      r_out(102)<=(mode and fifo_out(102)) or ((not mode) and ('0' xor fifo_out(11) xor fifo_out(102) xor fifo_out(120) xor fifo_out(180) xor fifo_out(229)));
      r_out(103)<=(mode and fifo_out(103)) or ((not mode) and ('0' xor fifo_out(233) xor fifo_out(27) xor fifo_out(45) xor fifo_out(103) xor fifo_out(217)));
      r_out(104)<=(mode and fifo_out(104)) or ((not mode) and ('0' xor fifo_out(8) xor fifo_out(44) xor fifo_out(104) xor fifo_out(124) xor fifo_out(135)));
      r_out(105)<=(mode and fifo_out(105)) or ((not mode) and ('0' xor fifo_out(75) xor fifo_out(100) xor fifo_out(105) xor fifo_out(161) xor fifo_out(172)));
      r_out(106)<=(mode and fifo_out(106)) or ((not mode) and ('0' xor fifo_out(57) xor fifo_out(91) xor fifo_out(106) xor fifo_out(187) xor fifo_out(194)));
      r_out(107)<=(mode and fifo_out(107)) or ((not mode) and ('0' xor fifo_out(73) xor fifo_out(93) xor fifo_out(107) xor fifo_out(156) xor fifo_out(198)));
      r_out(108)<=(mode and fifo_out(108)) or ((not mode) and ('0' xor fifo_out(0) xor fifo_out(28) xor fifo_out(99) xor fifo_out(108) xor fifo_out(190)));
      r_out(109)<=(mode and fifo_out(109)) or ((not mode) and ('0' xor fifo_out(40) xor fifo_out(51) xor fifo_out(109) xor fifo_out(193) xor fifo_out(205)));
      r_out(110)<=(mode and fifo_out(110)) or ((not mode) and ('0' xor fifo_out(27) xor fifo_out(67) xor fifo_out(110) xor fifo_out(162) xor fifo_out(177)));
      r_out(111)<=(mode and fifo_out(111)) or ((not mode) and ('0' xor fifo_out(47) xor fifo_out(60) xor fifo_out(71) xor fifo_out(111) xor fifo_out(231)));
      r_out(112)<=(mode and fifo_out(112)) or ((not mode) and ('0' xor fifo_out(31) xor fifo_out(105) xor fifo_out(112) xor fifo_out(119) xor fifo_out(219)));
      r_out(113)<=(mode and fifo_out(113)) or ((not mode) and ('0' xor fifo_out(89) xor fifo_out(95) xor fifo_out(113) xor fifo_out(118) xor fifo_out(127)));
      r_out(114)<=(mode and fifo_out(114)) or ((not mode) and ('0' xor fifo_out(24) xor fifo_out(59) xor fifo_out(114) xor fifo_out(157) xor fifo_out(195)));
      r_out(115)<=(mode and fifo_out(115)) or ((not mode) and ('0' xor fifo_out(42) xor fifo_out(92) xor fifo_out(115) xor fifo_out(117) xor fifo_out(189)));
      r_out(116)<=(mode and fifo_out(116)) or ((not mode) and ('0' xor fifo_out(116) xor fifo_out(162) xor fifo_out(184) xor fifo_out(191) xor fifo_out(224)));
      r_out(117)<=(mode and fifo_out(117)) or ((not mode) and ('0' xor fifo_out(42) xor fifo_out(72) xor fifo_out(77) xor fifo_out(117) xor fifo_out(182)));
      r_out(118)<=(mode and fifo_out(118)) or ((not mode) and ('0' xor fifo_out(53) xor fifo_out(95) xor fifo_out(118) xor fifo_out(200) xor fifo_out(227)));
      r_out(119)<=(mode and fifo_out(119)) or ((not mode) and ('0' xor fifo_out(18) xor fifo_out(119) xor fifo_out(147) xor fifo_out(158) xor fifo_out(166)));
      r_out(120)<=(mode and fifo_out(120)) or ((not mode) and ('0' xor fifo_out(24) xor fifo_out(25) xor fifo_out(120) xor fifo_out(180) xor fifo_out(195)));
      r_out(121)<=(mode and fifo_out(121)) or ((not mode) and ('0' xor fifo_out(106) xor fifo_out(119) xor fifo_out(121) xor fifo_out(144) xor fifo_out(179)));
      r_out(122)<=(mode and fifo_out(122)) or ((not mode) and ('0' xor fifo_out(48) xor fifo_out(76) xor fifo_out(107) xor fifo_out(122) xor fifo_out(145)));
      r_out(123)<=(mode and fifo_out(123)) or ((not mode) and ('0' xor fifo_out(16) xor fifo_out(86) xor fifo_out(94) xor fifo_out(123) xor fifo_out(128)));
      r_out(124)<=(mode and fifo_out(124)) or ((not mode) and ('0' xor fifo_out(12) xor fifo_out(31) xor fifo_out(124) xor fifo_out(140) xor fifo_out(151)));
      r_out(125)<=(mode and fifo_out(125)) or ((not mode) and ('0' xor fifo_out(69) xor fifo_out(120) xor fifo_out(125) xor fifo_out(133) xor fifo_out(198)));
      r_out(126)<=(mode and fifo_out(126)) or ((not mode) and ('0' xor fifo_out(19) xor fifo_out(42) xor fifo_out(81) xor fifo_out(121) xor fifo_out(126)));
      r_out(127)<=(mode and fifo_out(127)) or ((not mode) and ('0' xor fifo_out(14) xor fifo_out(49) xor fifo_out(50) xor fifo_out(127) xor fifo_out(173)));
      r_out(128)<=(mode and fifo_out(128)) or ((not mode) and ('0' xor fifo_out(7) xor fifo_out(98) xor fifo_out(128) xor fifo_out(150) xor fifo_out(161)));
      r_out(129)<=(mode and fifo_out(129)) or ((not mode) and ('0' xor fifo_out(8) xor fifo_out(60) xor fifo_out(89) xor fifo_out(122) xor fifo_out(129)));
      r_out(130)<=(mode and fifo_out(130)) or ((not mode) and ('0' xor fifo_out(10) xor fifo_out(90) xor fifo_out(130) xor fifo_out(137) xor fifo_out(175)));
      r_out(131)<=(mode and fifo_out(131)) or ((not mode) and ('0' xor fifo_out(121) xor fifo_out(131) xor fifo_out(135) xor fifo_out(156) xor fifo_out(199)));
      r_out(132)<=(mode and fifo_out(132)) or ((not mode) and ('0' xor fifo_out(41) xor fifo_out(93) xor fifo_out(110) xor fifo_out(132) xor fifo_out(231)));
      r_out(133)<=(mode and fifo_out(133)) or ((not mode) and ('0' xor fifo_out(4) xor fifo_out(6) xor fifo_out(43) xor fifo_out(133) xor fifo_out(165)));
      r_out(134)<=(mode and fifo_out(134)) or ((not mode) and ('0' xor fifo_out(2) xor fifo_out(53) xor fifo_out(72) xor fifo_out(82) xor fifo_out(134)));
      r_out(135)<=(mode and fifo_out(135)) or ((not mode) and ('0' xor fifo_out(56) xor fifo_out(104) xor fifo_out(135) xor fifo_out(143) xor fifo_out(190)));
      r_out(136)<=(mode and fifo_out(136)) or ((not mode) and ('0' xor fifo_out(5) xor fifo_out(127) xor fifo_out(136) xor fifo_out(140) xor fifo_out(208)));
      r_out(137)<=(mode and fifo_out(137)) or ((not mode) and ('0' xor fifo_out(37) xor fifo_out(68) xor fifo_out(137) xor fifo_out(159) xor fifo_out(214)));
      r_out(138)<=(mode and fifo_out(138)) or ((not mode) and ('0' xor fifo_out(82) xor fifo_out(92) xor fifo_out(104) xor fifo_out(138) xor fifo_out(145)));
      r_out(139)<=(mode and fifo_out(139)) or ((not mode) and ('0' xor fifo_out(29) xor fifo_out(36) xor fifo_out(83) xor fifo_out(139) xor fifo_out(181)));
      r_out(140)<=(mode and fifo_out(140)) or ((not mode) and ('0' xor fifo_out(12) xor fifo_out(95) xor fifo_out(140) xor fifo_out(168)));
      r_out(141)<=(mode and fifo_out(141)) or ((not mode) and ('0' xor fifo_out(233) xor fifo_out(141) xor fifo_out(156) xor fifo_out(183) xor fifo_out(186)));
      r_out(142)<=(mode and fifo_out(142)) or ((not mode) and ('0' xor fifo_out(26) xor fifo_out(108) xor fifo_out(142) xor fifo_out(163) xor fifo_out(173)));
      r_out(143)<=(mode and fifo_out(143)) or ((not mode) and ('0' xor fifo_out(52) xor fifo_out(103) xor fifo_out(139) xor fifo_out(143) xor fifo_out(147)));
      r_out(144)<=(mode and fifo_out(144)) or ((not mode) and ('0' xor fifo_out(1) xor fifo_out(125) xor fifo_out(144) xor fifo_out(218) xor fifo_out(223)));
      r_out(145)<=(mode and fifo_out(145)) or ((not mode) and ('0' xor fifo_out(37) xor fifo_out(75) xor fifo_out(145) xor fifo_out(176) xor fifo_out(188)));
      r_out(146)<=(mode and fifo_out(146)) or ((not mode) and ('0' xor fifo_out(43) xor fifo_out(133) xor fifo_out(146) xor fifo_out(175) xor fifo_out(188)));
      r_out(147)<=(mode and fifo_out(147)) or ((not mode) and ('0' xor fifo_out(87) xor fifo_out(147) xor fifo_out(154) xor fifo_out(168) xor fifo_out(223)));
      r_out(148)<=(mode and fifo_out(148)) or ((not mode) and ('0' xor fifo_out(19) xor fifo_out(41) xor fifo_out(49) xor fifo_out(123) xor fifo_out(148)));
      r_out(149)<=(mode and fifo_out(149)) or ((not mode) and ('0' xor fifo_out(106) xor fifo_out(141) xor fifo_out(143) xor fifo_out(149) xor fifo_out(179)));
      r_out(150)<=(mode and fifo_out(150)) or ((not mode) and ('0' xor fifo_out(68) xor fifo_out(87) xor fifo_out(136) xor fifo_out(150) xor fifo_out(177)));
      r_out(151)<=(mode and fifo_out(151)) or ((not mode) and ('0' xor fifo_out(101) xor fifo_out(151) xor fifo_out(167) xor fifo_out(223) xor fifo_out(227)));
      r_out(152)<=(mode and fifo_out(152)) or ((not mode) and ('0' xor fifo_out(20) xor fifo_out(32) xor fifo_out(76) xor fifo_out(152) xor fifo_out(230)));
      r_out(153)<=(mode and fifo_out(153)) or ((not mode) and ('0' xor fifo_out(100) xor fifo_out(137) xor fifo_out(153) xor fifo_out(171) xor fifo_out(190)));
      r_out(154)<=(mode and fifo_out(154)) or ((not mode) and ('0' xor fifo_out(14) xor fifo_out(71) xor fifo_out(114) xor fifo_out(154) xor fifo_out(195)));
      r_out(155)<=(mode and fifo_out(155)) or ((not mode) and ('0' xor fifo_out(65) xor fifo_out(123) xor fifo_out(155) xor fifo_out(178) xor fifo_out(196)));
      r_out(156)<=(mode and fifo_out(156)) or ((not mode) and ('0' xor fifo_out(233) xor fifo_out(64) xor fifo_out(131) xor fifo_out(156) xor fifo_out(229)));
      r_out(157)<=(mode and fifo_out(157)) or ((not mode) and ('0' xor fifo_out(95) xor fifo_out(109) xor fifo_out(152) xor fifo_out(157) xor fifo_out(170)));
      r_out(158)<=(mode and fifo_out(158)) or ((not mode) and ('0' xor fifo_out(100) xor fifo_out(113) xor fifo_out(134) xor fifo_out(158) xor fifo_out(214)));
      r_out(159)<=(mode and fifo_out(159)) or ((not mode) and ('0' xor fifo_out(29) xor fifo_out(64) xor fifo_out(159) xor fifo_out(187)));
      r_out(160)<=(mode and fifo_out(160)) or ((not mode) and ('0' xor fifo_out(33) xor fifo_out(65) xor fifo_out(90) xor fifo_out(119) xor fifo_out(160)));
      r_out(161)<=(mode and fifo_out(161)) or ((not mode) and ('0' xor fifo_out(118) xor fifo_out(161) xor fifo_out(170) xor fifo_out(178) xor fifo_out(197)));
      r_out(162)<=(mode and fifo_out(162)) or ((not mode) and ('0' xor fifo_out(19) xor fifo_out(75) xor fifo_out(147) xor fifo_out(162) xor fifo_out(207)));
      r_out(163)<=(mode and fifo_out(163)) or ((not mode) and ('0' xor fifo_out(114) xor fifo_out(115) xor fifo_out(163) xor fifo_out(184) xor fifo_out(216)));
      r_out(164)<=(mode and fifo_out(164)) or ((not mode) and ('0' xor fifo_out(7) xor fifo_out(56) xor fifo_out(88) xor fifo_out(148) xor fifo_out(164)));
      r_out(165)<=(mode and fifo_out(165)) or ((not mode) and ('0' xor fifo_out(143) xor fifo_out(165) xor fifo_out(181) xor fifo_out(193) xor fifo_out(204)));
      r_out(166)<=(mode and fifo_out(166)) or ((not mode) and ('0' xor fifo_out(54) xor fifo_out(89) xor fifo_out(92) xor fifo_out(162) xor fifo_out(166)));
      r_out(167)<=(mode and fifo_out(167)) or ((not mode) and ('0' xor fifo_out(5) xor fifo_out(52) xor fifo_out(61) xor fifo_out(167) xor fifo_out(174)));
      r_out(168)<=(mode and fifo_out(168)) or ((not mode) and ('0' xor fifo_out(14) xor fifo_out(41) xor fifo_out(119) xor fifo_out(168) xor fifo_out(179)));
      r_out(169)<=(mode and fifo_out(169)) or ((not mode) and ('0' xor fifo_out(26) xor fifo_out(36) xor fifo_out(117) xor fifo_out(169) xor fifo_out(216)));
      r_out(170)<=(mode and fifo_out(170)) or ((not mode) and ('0' xor fifo_out(66) xor fifo_out(170) xor fifo_out(172) xor fifo_out(181) xor fifo_out(206)));
      r_out(171)<=(mode and fifo_out(171)) or ((not mode) and ('0' xor fifo_out(118) xor fifo_out(125) xor fifo_out(139) xor fifo_out(155) xor fifo_out(171)));
      r_out(172)<=(mode and fifo_out(172)) or ((not mode) and ('0' xor fifo_out(8) xor fifo_out(30) xor fifo_out(127) xor fifo_out(142) xor fifo_out(172)));
      r_out(173)<=(mode and fifo_out(173)) or ((not mode) and ('0' xor fifo_out(61) xor fifo_out(78) xor fifo_out(173) xor fifo_out(209) xor fifo_out(232)));
      r_out(174)<=(mode and fifo_out(174)) or ((not mode) and ('0' xor fifo_out(34) xor fifo_out(98) xor fifo_out(112) xor fifo_out(133) xor fifo_out(174)));
      r_out(175)<=(mode and fifo_out(175)) or ((not mode) and ('0' xor fifo_out(4) xor fifo_out(102) xor fifo_out(160) xor fifo_out(175) xor fifo_out(212)));
      r_out(176)<=(mode and fifo_out(176)) or ((not mode) and ('0' xor fifo_out(125) xor fifo_out(160) xor fifo_out(176) xor fifo_out(195) xor fifo_out(209)));
      r_out(177)<=(mode and fifo_out(177)) or ((not mode) and ('0' xor fifo_out(63) xor fifo_out(105) xor fifo_out(136) xor fifo_out(177) xor fifo_out(208)));
      r_out(178)<=(mode and fifo_out(178)) or ((not mode) and ('0' xor fifo_out(39) xor fifo_out(73) xor fifo_out(129) xor fifo_out(163) xor fifo_out(178)));
      r_out(179)<=(mode and fifo_out(179)) or ((not mode) and ('0' xor fifo_out(66) xor fifo_out(102) xor fifo_out(118) xor fifo_out(179) xor fifo_out(182)));
      r_out(180)<=(mode and fifo_out(180)) or ((not mode) and ('0' xor fifo_out(20) xor fifo_out(139) xor fifo_out(151) xor fifo_out(176) xor fifo_out(180)));
      r_out(181)<=(mode and fifo_out(181)) or ((not mode) and ('0' xor fifo_out(2) xor fifo_out(5) xor fifo_out(70) xor fifo_out(151) xor fifo_out(181)));
      r_out(182)<=(mode and fifo_out(182)) or ((not mode) and ('0' xor fifo_out(17) xor fifo_out(22) xor fifo_out(69) xor fifo_out(138) xor fifo_out(182)));
      r_out(183)<=(mode and fifo_out(183)) or ((not mode) and ('0' xor fifo_out(2) xor fifo_out(20) xor fifo_out(40) xor fifo_out(55) xor fifo_out(183)));
      r_out(184)<=(mode and fifo_out(184)) or ((not mode) and ('0' xor fifo_out(10) xor fifo_out(49) xor fifo_out(70) xor fifo_out(94) xor fifo_out(184)));
      r_out(185)<=(mode and fifo_out(185)) or ((not mode) and ('0' xor fifo_out(96) xor fifo_out(103) xor fifo_out(174) xor fifo_out(185) xor fifo_out(222)));
      r_out(186)<=(mode and fifo_out(186)) or ((not mode) and ('0' xor fifo_out(21) xor fifo_out(63) xor fifo_out(85) xor fifo_out(186)));
      r_out(187)<=(mode and fifo_out(187)) or ((not mode) and ('0' xor fifo_out(16) xor fifo_out(53) xor fifo_out(91) xor fifo_out(160) xor fifo_out(187)));
      r_out(188)<=(mode and fifo_out(188)) or ((not mode) and ('0' xor fifo_out(1) xor fifo_out(35) xor fifo_out(53) xor fifo_out(149) xor fifo_out(188)));
      r_out(189)<=(mode and fifo_out(189)) or ((not mode) and ('0' xor fifo_out(0) xor fifo_out(33) xor fifo_out(189) xor fifo_out(200) xor fifo_out(211)));
      r_out(190)<=(mode and fifo_out(190)) or ((not mode) and ('0' xor fifo_out(7) xor fifo_out(98) xor fifo_out(131) xor fifo_out(190) xor fifo_out(203)));
      r_out(191)<=(mode and fifo_out(191)) or ((not mode) and ('0' xor fifo_out(1) xor fifo_out(34) xor fifo_out(87) xor fifo_out(115) xor fifo_out(191)));
      r_out(192)<=(mode and fifo_out(192)) or ((not mode) and ('0' xor fifo_out(30) xor fifo_out(59) xor fifo_out(167) xor fifo_out(187) xor fifo_out(192)));
      r_out(193)<=(mode and fifo_out(193)) or ((not mode) and ('0' xor fifo_out(30) xor fifo_out(78) xor fifo_out(103) xor fifo_out(193) xor fifo_out(220)));
      r_out(194)<=(mode and fifo_out(194)) or ((not mode) and ('0' xor fifo_out(135) xor fifo_out(179) xor fifo_out(185) xor fifo_out(187) xor fifo_out(194)));
      r_out(195)<=(mode and fifo_out(195)) or ((not mode) and ('0' xor fifo_out(55) xor fifo_out(109) xor fifo_out(112) xor fifo_out(195) xor fifo_out(215)));
      r_out(196)<=(mode and fifo_out(196)) or ((not mode) and ('0' xor fifo_out(80) xor fifo_out(97) xor fifo_out(182) xor fifo_out(196) xor fifo_out(210)));
      r_out(197)<=(mode and fifo_out(197)) or ((not mode) and ('0' xor fifo_out(12) xor fifo_out(105) xor fifo_out(117) xor fifo_out(197) xor fifo_out(214)));
      r_out(198)<=(mode and fifo_out(198)) or ((not mode) and ('0' xor fifo_out(100) xor fifo_out(104) xor fifo_out(129) xor fifo_out(198) xor fifo_out(205)));
      r_out(199)<=(mode and fifo_out(199)) or ((not mode) and ('0' xor fifo_out(2) xor fifo_out(84) xor fifo_out(124) xor fifo_out(163) xor fifo_out(199)));
      r_out(200)<=(mode and fifo_out(200)) or ((not mode) and ('0' xor fifo_out(56) xor fifo_out(85) xor fifo_out(126) xor fifo_out(200) xor fifo_out(230)));
      r_out(201)<=(mode and fifo_out(201)) or ((not mode) and ('0' xor fifo_out(104) xor fifo_out(150) xor fifo_out(180) xor fifo_out(201) xor fifo_out(212)));
      r_out(202)<=(mode and fifo_out(202)) or ((not mode) and ('0' xor fifo_out(13) xor fifo_out(76) xor fifo_out(79) xor fifo_out(202) xor fifo_out(231)));
      r_out(203)<=(mode and fifo_out(203)) or ((not mode) and ('0' xor fifo_out(28) xor fifo_out(51) xor fifo_out(122) xor fifo_out(192) xor fifo_out(203)));
      r_out(204)<=(mode and fifo_out(204)) or ((not mode) and ('0' xor fifo_out(37) xor fifo_out(44) xor fifo_out(127) xor fifo_out(204)));
      r_out(205)<=(mode and fifo_out(205)) or ((not mode) and ('0' xor fifo_out(25) xor fifo_out(115) xor fifo_out(173) xor fifo_out(205) xor fifo_out(221)));
      r_out(206)<=(mode and fifo_out(206)) or ((not mode) and ('0' xor fifo_out(23) xor fifo_out(201) xor fifo_out(203) xor fifo_out(206) xor fifo_out(224)));
      r_out(207)<=(mode and fifo_out(207)) or ((not mode) and ('0' xor fifo_out(14) xor fifo_out(73) xor fifo_out(149) xor fifo_out(163) xor fifo_out(207)));
      r_out(208)<=(mode and fifo_out(208)) or ((not mode) and ('0' xor fifo_out(106) xor fifo_out(166) xor fifo_out(197) xor fifo_out(208) xor fifo_out(225)));
      r_out(209)<=(mode and fifo_out(209)) or ((not mode) and ('0' xor fifo_out(44) xor fifo_out(66) xor fifo_out(125) xor fifo_out(170) xor fifo_out(209)));
      r_out(210)<=(mode and fifo_out(210)) or ((not mode) and ('0' xor fifo_out(45) xor fifo_out(63) xor fifo_out(101) xor fifo_out(210) xor fifo_out(228)));
      r_out(211)<=(mode and fifo_out(211)) or ((not mode) and ('0' xor fifo_out(29) xor fifo_out(47) xor fifo_out(149) xor fifo_out(201) xor fifo_out(211)));
      r_out(212)<=(mode and fifo_out(212)) or ((not mode) and ('0' xor fifo_out(68) xor fifo_out(148) xor fifo_out(174) xor fifo_out(212) xor fifo_out(215)));
      r_out(213)<=(mode and fifo_out(213)) or ((not mode) and ('0' xor fifo_out(18) xor fifo_out(178) xor fifo_out(193) xor fifo_out(213) xor fifo_out(228)));
      r_out(214)<=(mode and fifo_out(214)) or ((not mode) and ('0' xor fifo_out(55) xor fifo_out(158) xor fifo_out(183) xor fifo_out(214) xor fifo_out(222)));
      r_out(215)<=(mode and fifo_out(215)) or ((not mode) and ('0' xor fifo_out(43) xor fifo_out(46) xor fifo_out(111) xor fifo_out(114) xor fifo_out(215)));
      r_out(216)<=(mode and fifo_out(216)) or ((not mode) and ('0' xor fifo_out(0) xor fifo_out(46) xor fifo_out(216) xor fifo_out(217) xor fifo_out(229)));
      r_out(217)<=(mode and fifo_out(217)) or ((not mode) and ('0' xor fifo_out(15) xor fifo_out(19) xor fifo_out(37) xor fifo_out(216) xor fifo_out(217)));
      r_out(218)<=(mode and fifo_out(218)) or ((not mode) and ('0' xor fifo_out(0) xor fifo_out(35) xor fifo_out(177) xor fifo_out(218) xor fifo_out(220)));
      r_out(219)<=(mode and fifo_out(219)) or ((not mode) and ('0' xor fifo_out(96) xor fifo_out(114) xor fifo_out(134) xor fifo_out(157) xor fifo_out(219)));
      r_out(220)<=(mode and fifo_out(220)) or ((not mode) and ('0' xor fifo_out(38) xor fifo_out(74) xor fifo_out(110) xor fifo_out(112) xor fifo_out(220)));
      r_out(221)<=(mode and fifo_out(221)) or ((not mode) and ('0' xor fifo_out(48) xor fifo_out(72) xor fifo_out(109) xor fifo_out(169) xor fifo_out(221)));
      r_out(222)<=(mode and fifo_out(222)) or ((not mode) and ('0' xor fifo_out(87) xor fifo_out(107) xor fifo_out(144) xor fifo_out(213) xor fifo_out(222)));
      r_out(223)<=(mode and fifo_out(223)) or ((not mode) and ('0' xor fifo_out(45) xor fifo_out(90) xor fifo_out(92) xor fifo_out(150) xor fifo_out(223)));
      r_out(224)<=(mode and fifo_out(224)) or ((not mode) and ('0' xor fifo_out(20) xor fifo_out(135) xor fifo_out(138) xor fifo_out(186) xor fifo_out(224)));
      r_out(225)<=(mode and fifo_out(225)) or ((not mode) and ('0' xor fifo_out(111) xor fifo_out(202) xor fifo_out(224) xor fifo_out(225) xor fifo_out(230)));
      r_out(226)<=(mode and fifo_out(226)) or ((not mode) and ('0' xor fifo_out(79) xor fifo_out(86) xor fifo_out(107) xor fifo_out(142) xor fifo_out(226)));
      r_out(227)<=(mode and fifo_out(227)) or ((not mode) and ('0' xor fifo_out(98) xor fifo_out(142) xor fifo_out(153) xor fifo_out(161) xor fifo_out(227)));
      r_out(228)<=(mode and fifo_out(228)) or ((not mode) and ('0' xor fifo_out(165) xor fifo_out(196) xor fifo_out(210) xor fifo_out(228)));
      r_out(229)<=(mode and fifo_out(229)) or ((not mode) and ('0' xor fifo_out(4) xor fifo_out(65) xor fifo_out(67) xor fifo_out(140) xor fifo_out(229)));
      r_out(230)<=(mode and fifo_out(230)) or ((not mode) and ('0' xor fifo_out(62) xor fifo_out(69) xor fifo_out(101) xor fifo_out(202) xor fifo_out(230)));
      r_out(231)<=(mode and fifo_out(231)) or ((not mode) and ('0' xor fifo_out(18) xor fifo_out(88) xor fifo_out(132) xor fifo_out(164) xor fifo_out(231)));
      r_out(232)<=(mode and fifo_out(232)) or ((not mode) and ('0' xor fifo_out(144) xor fifo_out(159) xor fifo_out(170) xor fifo_out(213) xor fifo_out(232)));
      r_out(233)<=(mode and fifo_out(233)) or ((not mode) and ('0' xor fifo_out(233) xor fifo_out(46) xor fifo_out(91) xor fifo_out(172) xor fifo_out(175)));
    end if; end if;
  end process;
  fifo_out(0) <= r_out(1);
  fifo_out(1) <= r_out(2);
  fifo_out(2) <= r_out(3);
  fifo_out(3) <= r_out(4);
  fifo_out(4) <= r_out(5);
  fifo_out(5) <= r_out(6);
  fifo_out(6) <= r_out(7);
  fifo_out(7) <= r_out(8);
  fifo_out(8) <= r_out(9);
  fifo_out(9) <= r_out(10);
  fifo_out(10) <= r_out(11);
  fifo_out(11) <= r_out(12);
  fifo_out(12) <= r_out(13);
  fifo_out(13) <= r_out(14);
  fifo_out(14) <= r_out(15);
  fifo_out(15) <= r_out(16);
  fifo_out(16) <= r_out(17);
  fifo_out(17) <= r_out(18);
  fifo_out(18) <= r_out(19);
  fifo_out(19) <= r_out(20);
  fifo_out(20) <= r_out(21);
  fifo_out(21) <= r_out(22);
  fifo_out(22) <= r_out(23);
  fifo_out(23) <= r_out(24);
  fifo_out(24) <= r_out(25);
  fifo_out(25) <= r_out(26);
  fifo_out(26) <= r_out(27);
  fifo_out(27) <= r_out(28);
  fifo_out(28) <= r_out(29);
  fifo_out(29) <= r_out(30);
  fifo_out(30) <= r_out(31);
  fifo_out(31) <= r_out(32);
  fifo_out(32) <= r_out(33);
  fifo_out(33) <= r_out(34);
  fifo_out(34) <= r_out(35);
  fifo_out(35) <= r_out(36);
  fifo_out(36) <= r_out(37);
  fifo_out(37) <= r_out(38);
  fifo_out(38) <= r_out(39);
  fifo_out(39) <= r_out(40);
  fifo_out(40) <= r_out(41);
  fifo_out(41) <= r_out(42);
  fifo_out(42) <= r_out(43);
  fifo_out(43) <= r_out(44);
  fifo_out(44) <= r_out(45);
  fifo_out(45) <= r_out(46);
  fifo_out(46) <= r_out(47);
  fifo_out(47) <= r_out(48);
  fifo_out(48) <= r_out(49);
  fifo_out(49) <= r_out(50);
  fifo_out(50) <= r_out(51);
  fifo_out(51) <= r_out(52);
  fifo_out(52) <= r_out(53);
  fifo_out(53) <= r_out(54);
  fifo_out(54) <= r_out(55);
  fifo_out(55) <= r_out(56);
  fifo_out(56) <= r_out(57);
  fifo_out(57) <= r_out(58);
  fifo_out(58) <= r_out(59);
  fifo_out(59) <= r_out(60);
  fifo_out(60) <= r_out(61);
  fifo_out(61) <= r_out(62);
  fifo_out(62) <= r_out(63);
  fifo_out(63) <= r_out(64);
  fifo_out(64) <= r_out(65);
  fifo_out(65) <= r_out(66);
  fifo_out(66) <= r_out(67);
  fifo_out(67) <= r_out(68);
  fifo_out(68) <= r_out(69);
  fifo_out(69) <= r_out(70);
  fifo_out(70) <= r_out(71);
  fifo_out(71) <= r_out(72);
  fifo_out(72) <= r_out(73);
  fifo_out(73) <= r_out(74);
  fifo_out(74) <= r_out(75);
  fifo_out(75) <= r_out(76);
  fifo_out(76) <= r_out(77);
  fifo_out(77) <= r_out(78);
  fifo_out(78) <= r_out(79);
  fifo_out(79) <= r_out(80);
  fifo_out(80) <= r_out(81);
  fifo_out(81) <= r_out(82);
  fifo_out(82) <= r_out(83);
  fifo_out(83) <= r_out(84);
  fifo_out(84) <= r_out(85);
  fifo_out(85) <= r_out(86);
  fifo_out(86) <= r_out(87);
  fifo_out(87) <= r_out(88);
  fifo_out(88) <= r_out(89);
  fifo_out(89) <= r_out(90);
  fifo_out(90) <= r_out(91);
  fifo_out(91) <= r_out(92);
  fifo_out(92) <= r_out(93);
  fifo_out(93) <= r_out(94);
  fifo_out(94) <= r_out(95);
  fifo_out(95) <= r_out(96);
  fifo_out(96) <= r_out(97);
  fifo_out(97) <= r_out(98);
  fifo_out(98) <= r_out(99);
  fifo_out(99) <= r_out(100);
  fifo_out(100) <= r_out(101);
  fifo_out(101) <= r_out(102);
  fifo_out(102) <= r_out(103);
  fifo_out(103) <= r_out(104);
  fifo_out(104) <= r_out(105);
  fifo_out(105) <= r_out(106);
  fifo_out(106) <= r_out(107);
  fifo_out(107) <= r_out(108);
  fifo_out(108) <= r_out(109);
  fifo_out(109) <= r_out(110);
  fifo_out(110) <= r_out(111);
  fifo_out(111) <= r_out(112);
  fifo_out(112) <= r_out(113);
  fifo_out(113) <= r_out(114);
  fifo_out(114) <= r_out(115);
  fifo_out(115) <= r_out(116);
  fifo_out(116) <= r_out(117);
  fifo_out(117) <= r_out(118);
  fifo_out(118) <= r_out(119);
  fifo_out(119) <= r_out(120);
  fifo_out(120) <= r_out(121);
  fifo_out(121) <= r_out(122);
  fifo_out(122) <= r_out(123);
  fifo_out(123) <= r_out(124);
  fifo_out(124) <= r_out(125);
  fifo_out(125) <= r_out(126);
  fifo_out(126) <= r_out(127);
  fifo_out(127) <= r_out(128);
  fifo_out(128) <= r_out(129);
  fifo_out(129) <= r_out(130);
  fifo_out(130) <= r_out(131);
  fifo_out(131) <= r_out(132);
  fifo_out(132) <= r_out(133);
  fifo_out(133) <= r_out(134);
  fifo_out(134) <= r_out(135);
  fifo_out(135) <= r_out(136);
  fifo_out(136) <= r_out(137);
  fifo_out(137) <= r_out(138);
  fifo_out(138) <= r_out(139);
  fifo_out(139) <= r_out(140);
  fifo_out(140) <= r_out(141);
  fifo_out(141) <= r_out(142);
  fifo_out(142) <= r_out(143);
  fifo_out(143) <= r_out(144);
  fifo_out(144) <= r_out(145);
  fifo_out(145) <= r_out(146);
  fifo_out(146) <= r_out(147);
  fifo_out(147) <= r_out(148);
  fifo_out(148) <= r_out(149);
  fifo_out(149) <= r_out(150);
  fifo_out(150) <= r_out(151);
  fifo_out(151) <= r_out(152);
  fifo_out(152) <= r_out(153);
  fifo_out(153) <= r_out(154);
  fifo_out(154) <= r_out(155);
  fifo_out(155) <= r_out(156);
  fifo_out(156) <= r_out(157);
  fifo_out(157) <= r_out(158);
  fifo_out(158) <= r_out(159);
  fifo_out(159) <= r_out(160);
  fifo_out(160) <= r_out(161);
  fifo_out(161) <= r_out(162);
  fifo_out(162) <= r_out(163);
  fifo_out(163) <= r_out(164);
  fifo_out(164) <= r_out(165);
  fifo_out(165) <= r_out(166);
  fifo_out(166) <= r_out(167);
  fifo_out(167) <= r_out(168);
  fifo_out(168) <= r_out(169);
  fifo_out(169) <= r_out(170);
  fifo_out(170) <= r_out(171);
  fifo_out(171) <= r_out(172);
  fifo_out(172) <= r_out(173);
  fifo_out(173) <= r_out(174);
  fifo_out(174) <= r_out(175);
  fifo_out(175) <= r_out(176);
  fifo_out(176) <= r_out(177);
  fifo_out(177) <= r_out(178);
  fifo_out(178) <= r_out(179);
  fifo_out(179) <= r_out(180);
  fifo_out(180) <= r_out(181);
  fifo_out(181) <= r_out(182);
  fifo_out(182) <= r_out(183);
  fifo_out(183) <= r_out(184);
  fifo_out(184) <= r_out(185);
  fifo_out(185) <= r_out(186);
  fifo_out(186) <= r_out(187);
  fifo_out(187) <= r_out(188);
  fifo_out(188) <= r_out(189);
  fifo_out(189) <= r_out(190);
  fifo_out(190) <= r_out(191);
  fifo_out(191) <= r_out(192);
  fifo_out(192) <= r_out(193);
  fifo_out(193) <= r_out(194);
  fifo_out(194) <= r_out(195);
  fifo_out(195) <= r_out(196);
  fifo_out(196) <= r_out(197);
  fifo_out(197) <= r_out(198);
  fifo_out(198) <= r_out(199);
  fifo_out(199) <= r_out(200);
  fifo_out(200) <= r_out(201);
  fifo_out(201) <= r_out(202);
  fifo_out(202) <= r_out(203);
  fifo_out(203) <= r_out(204);
  fifo_out(204) <= r_out(205);
  fifo_out(205) <= r_out(206);
  fifo_out(206) <= r_out(207);
  fifo_out(207) <= r_out(208);
  fifo_out(208) <= r_out(209);
  fifo_out(209) <= r_out(210);
  fifo_out(210) <= r_out(211);
  fifo_out(211) <= r_out(212);
  fifo_out(212) <= r_out(213);
  fifo_out(213) <= r_out(214);
  fifo_out(214) <= r_out(215);
  fifo_out(215) <= r_out(216);
  fifo_out(216) <= r_out(217);
  fifo_out(217) <= r_out(218);
  fifo_out(218) <= r_out(219);
  fifo_out(219) <= r_out(220);
  fifo_out(220) <= r_out(221);
  fifo_out(221) <= r_out(222);
  fifo_out(222) <= r_out(223);
  fifo_out(223) <= r_out(224);
  fifo_out(224) <= r_out(225);
  fifo_out(225) <= r_out(226);
  fifo_out(226) <= r_out(227);
  fifo_out(227) <= r_out(228);
  fifo_out(228) <= r_out(229);
  fifo_out(229) <= r_out(230);
  fifo_out(230) <= r_out(231);
  fifo_out(231) <= r_out(232);
  fifo_out(232) <= r_out(233);
  fifo_out(233) <= r_out(0);
end RTL;
