
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;

package common is
constant LLR_BITS :natural := 6;
type llr_row_t is array(0 to 1-1) of signed(6-1 downto 0);
type llr_array_t is array(0 to 127-1, 0  to 1-1) of signed(6-1 downto 0);
type llr_column_t is array(0 to 127-1) of signed(6-1 downto 0);
subtype column_sum_t is signed(10-1 downto 0);
type column_sum_array_t is array(0 to 127-1) of column_sum_t;
subtype min_signs_t is std_logic_vector(0 to 127-1);
subtype min_t is unsigned(6-1 downto 0);
type min_array_t is array(0 to 127-1) of unsigned(6-1 downto 0);
type signs_t is array(0 to 127-1) of std_logic_vector(0 to 1-1);
subtype min_id_t is unsigned(5-1 downto 0);
type min_id_array_t is array(0 to 127-1) of min_id_t;
type roll_count_t is array(0 to 1-1) of natural;
subtype row_addr_t is unsigned(7-1 downto 0);
subtype col_addr_t is unsigned(6-1 downto 0);
subtype signs_addr_t is unsigned(9-1 downto 0);
subtype roll_t is unsigned(7-1 downto 0);
constant ROLL_COUNT : roll_count_t := (0, others => 0);
constant HQC_COLUMNS : natural := 66;
constant VN_MEM_BITS : natural := 7;
constant CN_MEM_BITS : natural := 6;
subtype vec_inst_t is std_logic_vector(80-1 downto 0);
type inst_t is 
    record
        row_end : std_logic;
        col_end : std_logic;
        llr_mem_rd : std_logic;
        llr_mem_addr : row_addr_t;
        result_addr : row_addr_t;
        result_wr : std_logic;
        store_cn_wr : std_logic;
        store_cn_addr : col_addr_t;
        load_cn_rd : std_logic;
        load_cn_addr : col_addr_t;
        store_vn_wr : std_logic;
        store_vn_addr : row_addr_t;
        load_vn_rd : std_logic;
        load_vn_addr : row_addr_t;
        store_signs_wr : std_logic;
        store_signs_addr : signs_addr_t;
        load_signs_rd : std_logic;
        load_signs_addr : signs_addr_t;
        min_offset : min_id_t;
        roll : roll_t;
    end record;
function pack(int_in : inst_t) return std_logic_vector;
function unpack(int_in : std_logic_vector) return inst_t;
type inst_array_t is array(integer range <>) of vec_inst_t;
constant INSTRUCTIONS : inst_array_t(0 to 704-1) := (pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000000000", min_offset => "00000", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000001", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000000001", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011010", store_signs_wr => '1',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000000010", min_offset => "00000", roll => "1100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011100", store_signs_wr => '1',store_signs_addr => "000000001", load_signs_rd => '1',load_signs_addr => "000000011", min_offset => "00001", roll => "1001101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100010", store_signs_wr => '1',store_signs_addr => "000000010", load_signs_rd => '1',load_signs_addr => "000000100", min_offset => "00010", roll => "1111011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001000", store_signs_wr => '1',store_signs_addr => "000000011", load_signs_rd => '1',load_signs_addr => "000000101", min_offset => "00011", roll => "1011100")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001010", store_signs_wr => '1',store_signs_addr => "000000100", load_signs_rd => '1',load_signs_addr => "000000110", min_offset => "00100", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001100", store_signs_wr => '1',store_signs_addr => "000000101", load_signs_rd => '1',load_signs_addr => "000000111", min_offset => "00000", roll => "0010110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001101", store_signs_wr => '1',store_signs_addr => "000000110", load_signs_rd => '1',load_signs_addr => "000001000", min_offset => "00001", roll => "1011010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011010", store_signs_wr => '1',store_signs_addr => "000000111", load_signs_rd => '1',load_signs_addr => "000001001", min_offset => "00010", roll => "1011110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100010", store_signs_wr => '1',store_signs_addr => "000001000", load_signs_rd => '1',load_signs_addr => "000001010", min_offset => "00011", roll => "0001000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100011", store_signs_wr => '1',store_signs_addr => "000001001", load_signs_rd => '1',load_signs_addr => "000001011", min_offset => "00100", roll => "0111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001000", store_signs_wr => '1',store_signs_addr => "000001010", load_signs_rd => '1',load_signs_addr => "000001100", min_offset => "00101", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "000001", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001101", store_signs_wr => '1',store_signs_addr => "000001011", load_signs_rd => '1',load_signs_addr => "000001101", min_offset => "00110", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011011", store_signs_wr => '1',store_signs_addr => "000001100", load_signs_rd => '1',load_signs_addr => "000001110", min_offset => "00000", roll => "1010111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011101", store_signs_wr => '1',store_signs_addr => "000001101", load_signs_rd => '1',load_signs_addr => "000001111", min_offset => "00001", roll => "0110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100011", store_signs_wr => '1',store_signs_addr => "000001110", load_signs_rd => '1',load_signs_addr => "000010000", min_offset => "00010", roll => "1010111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100100", store_signs_wr => '1',store_signs_addr => "000001111", load_signs_rd => '1',load_signs_addr => "000010001", min_offset => "00011", roll => "1110010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001111", store_signs_wr => '1',store_signs_addr => "000010000", load_signs_rd => '1',load_signs_addr => "000010010", min_offset => "00100", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "000010", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010011", store_signs_wr => '1',store_signs_addr => "000010001", load_signs_rd => '1',load_signs_addr => "000010011", min_offset => "00101", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011011", store_signs_wr => '1',store_signs_addr => "000010010", load_signs_rd => '1',load_signs_addr => "000010100", min_offset => "00000", roll => "1000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100000", store_signs_wr => '1',store_signs_addr => "000010011", load_signs_rd => '1',load_signs_addr => "000010101", min_offset => "00001", roll => "1000101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100100", store_signs_wr => '1',store_signs_addr => "000010100", load_signs_rd => '1',load_signs_addr => "000010110", min_offset => "00010", roll => "1111000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100101", store_signs_wr => '1',store_signs_addr => "000010101", load_signs_rd => '1',load_signs_addr => "000010111", min_offset => "00011", roll => "1101011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000111", store_signs_wr => '1',store_signs_addr => "000010110", load_signs_rd => '1',load_signs_addr => "000011000", min_offset => "00100", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "000011", load_cn_rd => '1',load_cn_addr => "000100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001000", store_signs_wr => '1',store_signs_addr => "000010111", load_signs_rd => '1',load_signs_addr => "000011001", min_offset => "00101", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010011", store_signs_wr => '1',store_signs_addr => "000011000", load_signs_rd => '1',load_signs_addr => "000011010", min_offset => "00000", roll => "1110000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100101", store_signs_wr => '1',store_signs_addr => "000011001", load_signs_rd => '1',load_signs_addr => "000011011", min_offset => "00001", roll => "1001111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100110", store_signs_wr => '1',store_signs_addr => "000011010", load_signs_rd => '1',load_signs_addr => "000011100", min_offset => "00010", roll => "1000011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001111", store_signs_wr => '1',store_signs_addr => "000011011", load_signs_rd => '1',load_signs_addr => "000011101", min_offset => "00011", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "000100", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010110", store_signs_wr => '1',store_signs_addr => "000011100", load_signs_rd => '1',load_signs_addr => "000011110", min_offset => "00100", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011010", store_signs_wr => '1',store_signs_addr => "000011101", load_signs_rd => '1',load_signs_addr => "000011111", min_offset => "00000", roll => "0111111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011011", store_signs_wr => '1',store_signs_addr => "000011110", load_signs_rd => '1',load_signs_addr => "000100000", min_offset => "00001", roll => "0111011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100110", store_signs_wr => '1',store_signs_addr => "000011111", load_signs_rd => '1',load_signs_addr => "000100001", min_offset => "00010", roll => "0101111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100111", store_signs_wr => '1',store_signs_addr => "000100000", load_signs_rd => '1',load_signs_addr => "000100010", min_offset => "00011", roll => "1000101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000001", store_signs_wr => '1',store_signs_addr => "000100001", load_signs_rd => '1',load_signs_addr => "000100011", min_offset => "00100", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "000101", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000011", store_signs_wr => '1',store_signs_addr => "000100010", load_signs_rd => '1',load_signs_addr => "000100100", min_offset => "00101", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000101", store_signs_wr => '1',store_signs_addr => "000100011", load_signs_rd => '1',load_signs_addr => "000100101", min_offset => "00000", roll => "1001100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001001", store_signs_wr => '1',store_signs_addr => "000100100", load_signs_rd => '1',load_signs_addr => "000100110", min_offset => "00001", roll => "0001110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001011", store_signs_wr => '1',store_signs_addr => "000100101", load_signs_rd => '1',load_signs_addr => "000100111", min_offset => "00010", roll => "0110001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001101", store_signs_wr => '1',store_signs_addr => "000100110", load_signs_rd => '1',load_signs_addr => "000101000", min_offset => "00011", roll => "1111000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010011", store_signs_wr => '1',store_signs_addr => "000100111", load_signs_rd => '1',load_signs_addr => "000101001", min_offset => "00100", roll => "1110110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011001", store_signs_wr => '1',store_signs_addr => "000101000", load_signs_rd => '1',load_signs_addr => "000101010", min_offset => "00101", roll => "1110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011101", store_signs_wr => '1',store_signs_addr => "000101001", load_signs_rd => '1',load_signs_addr => "000101011", min_offset => "00110", roll => "1100010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100000", store_signs_wr => '1',store_signs_addr => "000101010", load_signs_rd => '1',load_signs_addr => "000101100", min_offset => "00111", roll => "1111001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100110", store_signs_wr => '1',store_signs_addr => "000101011", load_signs_rd => '1',load_signs_addr => "000101101", min_offset => "01000", roll => "1001011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100111", store_signs_wr => '1',store_signs_addr => "000101100", load_signs_rd => '1',load_signs_addr => "000101110", min_offset => "01001", roll => "1101011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101000", store_signs_wr => '1',store_signs_addr => "000101101", load_signs_rd => '1',load_signs_addr => "000101111", min_offset => "01010", roll => "0000010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000101", store_signs_wr => '1',store_signs_addr => "000101110", load_signs_rd => '1',load_signs_addr => "000110000", min_offset => "01011", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "000110", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000111", store_signs_wr => '1',store_signs_addr => "000101111", load_signs_rd => '1',load_signs_addr => "000110001", min_offset => "01100", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001100", store_signs_wr => '1',store_signs_addr => "000110000", load_signs_rd => '1',load_signs_addr => "000110010", min_offset => "00000", roll => "0011111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001101", store_signs_wr => '1',store_signs_addr => "000110001", load_signs_rd => '1',load_signs_addr => "000110011", min_offset => "00001", roll => "0110010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010000", store_signs_wr => '1',store_signs_addr => "000110010", load_signs_rd => '1',load_signs_addr => "000110100", min_offset => "00010", roll => "0001111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010010", store_signs_wr => '1',store_signs_addr => "000110011", load_signs_rd => '1',load_signs_addr => "000110101", min_offset => "00011", roll => "0111111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010110", store_signs_wr => '1',store_signs_addr => "000110100", load_signs_rd => '1',load_signs_addr => "000110110", min_offset => "00100", roll => "0000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010111", store_signs_wr => '1',store_signs_addr => "000110101", load_signs_rd => '1',load_signs_addr => "000110111", min_offset => "00101", roll => "0000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100000", store_signs_wr => '1',store_signs_addr => "000110110", load_signs_rd => '1',load_signs_addr => "000111000", min_offset => "00110", roll => "1100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100010", store_signs_wr => '1',store_signs_addr => "000110111", load_signs_rd => '1',load_signs_addr => "000111001", min_offset => "00111", roll => "1100011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100110", store_signs_wr => '1',store_signs_addr => "000111000", load_signs_rd => '1',load_signs_addr => "000111010", min_offset => "01000", roll => "1100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101000", store_signs_wr => '1',store_signs_addr => "000111001", load_signs_rd => '1',load_signs_addr => "000111011", min_offset => "01001", roll => "1110001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101001", store_signs_wr => '1',store_signs_addr => "000111010", load_signs_rd => '1',load_signs_addr => "000111100", min_offset => "01010", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000010", store_signs_wr => '1',store_signs_addr => "000111011", load_signs_rd => '1',load_signs_addr => "000111101", min_offset => "01011", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "000111", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001011", store_signs_wr => '1',store_signs_addr => "000111100", load_signs_rd => '1',load_signs_addr => "000111110", min_offset => "01100", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001110", store_signs_wr => '1',store_signs_addr => "000111101", load_signs_rd => '1',load_signs_addr => "000111111", min_offset => "00000", roll => "1000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001111", store_signs_wr => '1',store_signs_addr => "000111110", load_signs_rd => '1',load_signs_addr => "001000000", min_offset => "00001", roll => "0101001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010011", store_signs_wr => '1',store_signs_addr => "000111111", load_signs_rd => '1',load_signs_addr => "001000001", min_offset => "00010", roll => "1001100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011001", store_signs_wr => '1',store_signs_addr => "001000000", load_signs_rd => '1',load_signs_addr => "001000010", min_offset => "00011", roll => "0101111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011010", store_signs_wr => '1',store_signs_addr => "001000001", load_signs_rd => '1',load_signs_addr => "001000011", min_offset => "00100", roll => "1101101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011011", store_signs_wr => '1',store_signs_addr => "001000010", load_signs_rd => '1',load_signs_addr => "001000100", min_offset => "00101", roll => "0111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011101", store_signs_wr => '1',store_signs_addr => "001000011", load_signs_rd => '1',load_signs_addr => "001000101", min_offset => "00110", roll => "1110000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101001", store_signs_wr => '1',store_signs_addr => "001000100", load_signs_rd => '1',load_signs_addr => "001000110", min_offset => "00111", roll => "1110100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101010", store_signs_wr => '1',store_signs_addr => "001000101", load_signs_rd => '1',load_signs_addr => "001000111", min_offset => "01000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000010", store_signs_wr => '1',store_signs_addr => "001000110", load_signs_rd => '1',load_signs_addr => "001001000", min_offset => "01001", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "001000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001010", store_signs_wr => '1',store_signs_addr => "001000111", load_signs_rd => '1',load_signs_addr => "001001001", min_offset => "01010", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001110", store_signs_wr => '1',store_signs_addr => "001001000", load_signs_rd => '1',load_signs_addr => "001001010", min_offset => "00000", roll => "0110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010001", store_signs_wr => '1',store_signs_addr => "001001001", load_signs_rd => '1',load_signs_addr => "001001011", min_offset => "00001", roll => "0111100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010010", store_signs_wr => '1',store_signs_addr => "001001010", load_signs_rd => '1',load_signs_addr => "001001100", min_offset => "00010", roll => "0101110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011001", store_signs_wr => '1',store_signs_addr => "001001011", load_signs_rd => '1',load_signs_addr => "001001101", min_offset => "00011", roll => "1001011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011011", store_signs_wr => '1',store_signs_addr => "001001100", load_signs_rd => '1',load_signs_addr => "001001110", min_offset => "00100", roll => "0100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011111", store_signs_wr => '1',store_signs_addr => "001001101", load_signs_rd => '1',load_signs_addr => "001001111", min_offset => "00101", roll => "0111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100101", store_signs_wr => '1',store_signs_addr => "001001110", load_signs_rd => '1',load_signs_addr => "001010000", min_offset => "00110", roll => "1010011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101001", store_signs_wr => '1',store_signs_addr => "001001111", load_signs_rd => '1',load_signs_addr => "001010001", min_offset => "00111", roll => "1101101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101010", store_signs_wr => '1',store_signs_addr => "001010000", load_signs_rd => '1',load_signs_addr => "001010010", min_offset => "01000", roll => "0110001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101011", store_signs_wr => '1',store_signs_addr => "001010001", load_signs_rd => '1',load_signs_addr => "001010011", min_offset => "01001", roll => "0110111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000000", store_signs_wr => '1',store_signs_addr => "001010010", load_signs_rd => '1',load_signs_addr => "001010100", min_offset => "01010", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "001001", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000001", store_signs_wr => '1',store_signs_addr => "001010011", load_signs_rd => '1',load_signs_addr => "001010101", min_offset => "01011", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000010", store_signs_wr => '1',store_signs_addr => "001010100", load_signs_rd => '1',load_signs_addr => "001010110", min_offset => "00000", roll => "0101010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001100", store_signs_wr => '1',store_signs_addr => "001010101", load_signs_rd => '1',load_signs_addr => "001010111", min_offset => "00001", roll => "1000010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011110", store_signs_wr => '1',store_signs_addr => "001010110", load_signs_rd => '1',load_signs_addr => "001011000", min_offset => "00010", roll => "1101111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011111", store_signs_wr => '1',store_signs_addr => "001010111", load_signs_rd => '1',load_signs_addr => "001011001", min_offset => "00011", roll => "0110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100111", store_signs_wr => '1',store_signs_addr => "001011000", load_signs_rd => '1',load_signs_addr => "001011010", min_offset => "00100", roll => "0101001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101011", store_signs_wr => '1',store_signs_addr => "001011001", load_signs_rd => '1',load_signs_addr => "001011011", min_offset => "00101", roll => "1110000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101100", store_signs_wr => '1',store_signs_addr => "001011010", load_signs_rd => '1',load_signs_addr => "001011100", min_offset => "00110", roll => "0101100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000111", store_signs_wr => '1',store_signs_addr => "001011011", load_signs_rd => '1',load_signs_addr => "001011101", min_offset => "00111", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "001010", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001101", store_signs_wr => '1',store_signs_addr => "001011100", load_signs_rd => '1',load_signs_addr => "001011110", min_offset => "01000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011001", store_signs_wr => '1',store_signs_addr => "001011101", load_signs_rd => '1',load_signs_addr => "001011111", min_offset => "00000", roll => "0000010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011010", store_signs_wr => '1',store_signs_addr => "001011110", load_signs_rd => '1',load_signs_addr => "001100000", min_offset => "00001", roll => "1101001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011110", store_signs_wr => '1',store_signs_addr => "001011111", load_signs_rd => '1',load_signs_addr => "001100001", min_offset => "00010", roll => "1111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011111", store_signs_wr => '1',store_signs_addr => "001100000", load_signs_rd => '1',load_signs_addr => "001100010", min_offset => "00011", roll => "1001001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100000", store_signs_wr => '1',store_signs_addr => "001100001", load_signs_rd => '1',load_signs_addr => "001100011", min_offset => "00100", roll => "1000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100100", store_signs_wr => '1',store_signs_addr => "001100010", load_signs_rd => '1',load_signs_addr => "001100100", min_offset => "00101", roll => "1010111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101100", store_signs_wr => '1',store_signs_addr => "001100011", load_signs_rd => '1',load_signs_addr => "001100101", min_offset => "00110", roll => "1100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101101", store_signs_wr => '1',store_signs_addr => "001100100", load_signs_rd => '1',load_signs_addr => "001100110", min_offset => "00111", roll => "0100001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001110", store_signs_wr => '1',store_signs_addr => "001100101", load_signs_rd => '1',load_signs_addr => "001100111", min_offset => "01000", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "001011", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010100", store_signs_wr => '1',store_signs_addr => "001100110", load_signs_rd => '1',load_signs_addr => "001101000", min_offset => "01001", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011011", store_signs_wr => '1',store_signs_addr => "001100111", load_signs_rd => '1',load_signs_addr => "001101001", min_offset => "00000", roll => "0110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100101", store_signs_wr => '1',store_signs_addr => "001101000", load_signs_rd => '1',load_signs_addr => "001101010", min_offset => "00001", roll => "1000011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100110", store_signs_wr => '1',store_signs_addr => "001101001", load_signs_rd => '1',load_signs_addr => "001101011", min_offset => "00010", roll => "1000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101100", store_signs_wr => '1',store_signs_addr => "001101010", load_signs_rd => '1',load_signs_addr => "001101100", min_offset => "00011", roll => "1110110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101101", store_signs_wr => '1',store_signs_addr => "001101011", load_signs_rd => '1',load_signs_addr => "001101101", min_offset => "00100", roll => "1111101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101110", store_signs_wr => '1',store_signs_addr => "001101100", load_signs_rd => '1',load_signs_addr => "001101110", min_offset => "00101", roll => "1001101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000010", store_signs_wr => '1',store_signs_addr => "001101101", load_signs_rd => '1',load_signs_addr => "001101111", min_offset => "00110", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "001100", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000110", store_signs_wr => '1',store_signs_addr => "001101110", load_signs_rd => '1',load_signs_addr => "001110000", min_offset => "00111", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000111", store_signs_wr => '1',store_signs_addr => "001101111", load_signs_rd => '1',load_signs_addr => "001110001", min_offset => "00000", roll => "1011001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001111", store_signs_wr => '1',store_signs_addr => "001110000", load_signs_rd => '1',load_signs_addr => "001110010", min_offset => "00001", roll => "1000101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100000", store_signs_wr => '1',store_signs_addr => "001110001", load_signs_rd => '1',load_signs_addr => "001110011", min_offset => "00010", roll => "1011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101001", store_signs_wr => '1',store_signs_addr => "001110010", load_signs_rd => '1',load_signs_addr => "001110100", min_offset => "00011", roll => "1011111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101110", store_signs_wr => '1',store_signs_addr => "001110011", load_signs_rd => '1',load_signs_addr => "001110101", min_offset => "00100", roll => "0101101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101111", store_signs_wr => '1',store_signs_addr => "001110100", load_signs_rd => '1',load_signs_addr => "001110110", min_offset => "00101", roll => "0111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000100", store_signs_wr => '1',store_signs_addr => "001110101", load_signs_rd => '1',load_signs_addr => "001110111", min_offset => "00110", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "001101", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000111", store_signs_wr => '1',store_signs_addr => "001110110", load_signs_rd => '1',load_signs_addr => "001111000", min_offset => "00111", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001010", store_signs_wr => '1',store_signs_addr => "001110111", load_signs_rd => '1',load_signs_addr => "001111001", min_offset => "00000", roll => "1100000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001101", store_signs_wr => '1',store_signs_addr => "001111000", load_signs_rd => '1',load_signs_addr => "001111010", min_offset => "00001", roll => "0111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010000", store_signs_wr => '1',store_signs_addr => "001111001", load_signs_rd => '1',load_signs_addr => "001111011", min_offset => "00010", roll => "0000110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010010", store_signs_wr => '1',store_signs_addr => "001111010", load_signs_rd => '1',load_signs_addr => "001111100", min_offset => "00011", roll => "1101111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010100", store_signs_wr => '1',store_signs_addr => "001111011", load_signs_rd => '1',load_signs_addr => "001111101", min_offset => "00100", roll => "0110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100011", store_signs_wr => '1',store_signs_addr => "001111100", load_signs_rd => '1',load_signs_addr => "001111110", min_offset => "00101", roll => "0100111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101111", store_signs_wr => '1',store_signs_addr => "001111101", load_signs_rd => '1',load_signs_addr => "001111111", min_offset => "00110", roll => "0111001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110000", store_signs_wr => '1',store_signs_addr => "001111110", load_signs_rd => '1',load_signs_addr => "010000000", min_offset => "00111", roll => "0010110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000010", store_signs_wr => '1',store_signs_addr => "001111111", load_signs_rd => '1',load_signs_addr => "010000001", min_offset => "01000", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "001110", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000101", store_signs_wr => '1',store_signs_addr => "010000000", load_signs_rd => '1',load_signs_addr => "010000010", min_offset => "01001", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001001", store_signs_wr => '1',store_signs_addr => "010000001", load_signs_rd => '1',load_signs_addr => "010000011", min_offset => "00000", roll => "1000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001100", store_signs_wr => '1',store_signs_addr => "010000010", load_signs_rd => '1',load_signs_addr => "010000100", min_offset => "00001", roll => "0001001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001110", store_signs_wr => '1',store_signs_addr => "010000011", load_signs_rd => '1',load_signs_addr => "010000101", min_offset => "00010", roll => "1000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010010", store_signs_wr => '1',store_signs_addr => "010000100", load_signs_rd => '1',load_signs_addr => "010000110", min_offset => "00011", roll => "1011011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010111", store_signs_wr => '1',store_signs_addr => "010000101", load_signs_rd => '1',load_signs_addr => "010000111", min_offset => "00100", roll => "0111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011000", store_signs_wr => '1',store_signs_addr => "010000110", load_signs_rd => '1',load_signs_addr => "010001000", min_offset => "00101", roll => "0010010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011001", store_signs_wr => '1',store_signs_addr => "010000111", load_signs_rd => '1',load_signs_addr => "010001001", min_offset => "00110", roll => "0100111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100000", store_signs_wr => '1',store_signs_addr => "010001000", load_signs_rd => '1',load_signs_addr => "010001010", min_offset => "00111", roll => "1000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100010", store_signs_wr => '1',store_signs_addr => "010001001", load_signs_rd => '1',load_signs_addr => "010001011", min_offset => "01000", roll => "0000100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100101", store_signs_wr => '1',store_signs_addr => "010001010", load_signs_rd => '1',load_signs_addr => "010001100", min_offset => "01001", roll => "0010100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110000", store_signs_wr => '1',store_signs_addr => "010001011", load_signs_rd => '1',load_signs_addr => "010001101", min_offset => "01010", roll => "1011110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110001", store_signs_wr => '1',store_signs_addr => "010001100", load_signs_rd => '1',load_signs_addr => "010001110", min_offset => "01011", roll => "1010011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001110", store_signs_wr => '1',store_signs_addr => "010001101", load_signs_rd => '1',load_signs_addr => "010001111", min_offset => "01100", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "001111", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011110", store_signs_wr => '1',store_signs_addr => "010001110", load_signs_rd => '1',load_signs_addr => "010010000", min_offset => "01101", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100111", store_signs_wr => '1',store_signs_addr => "010001111", load_signs_rd => '1',load_signs_addr => "010010001", min_offset => "00000", roll => "1110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110000", store_signs_wr => '1',store_signs_addr => "010010000", load_signs_rd => '1',load_signs_addr => "010010010", min_offset => "00001", roll => "1000010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110001", store_signs_wr => '1',store_signs_addr => "010010001", load_signs_rd => '1',load_signs_addr => "010010011", min_offset => "00010", roll => "0100100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110010", store_signs_wr => '1',store_signs_addr => "010010010", load_signs_rd => '1',load_signs_addr => "010010100", min_offset => "00011", roll => "0101011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000011", store_signs_wr => '1',store_signs_addr => "010010011", load_signs_rd => '1',load_signs_addr => "010010101", min_offset => "00100", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "010000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000100", store_signs_wr => '1',store_signs_addr => "010010100", load_signs_rd => '1',load_signs_addr => "010010110", min_offset => "00101", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000111", store_signs_wr => '1',store_signs_addr => "010010101", load_signs_rd => '1',load_signs_addr => "010010111", min_offset => "00000", roll => "0111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001000", store_signs_wr => '1',store_signs_addr => "010010110", load_signs_rd => '1',load_signs_addr => "010011000", min_offset => "00001", roll => "1110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010100", store_signs_wr => '1',store_signs_addr => "010010111", load_signs_rd => '1',load_signs_addr => "010011001", min_offset => "00010", roll => "0110110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010110", store_signs_wr => '1',store_signs_addr => "010011000", load_signs_rd => '1',load_signs_addr => "010011010", min_offset => "00011", roll => "0100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011011", store_signs_wr => '1',store_signs_addr => "010011001", load_signs_rd => '1',load_signs_addr => "010011011", min_offset => "00100", roll => "0100111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011101", store_signs_wr => '1',store_signs_addr => "010011010", load_signs_rd => '1',load_signs_addr => "010011100", min_offset => "00101", roll => "1011100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011110", store_signs_wr => '1',store_signs_addr => "010011011", load_signs_rd => '1',load_signs_addr => "010011101", min_offset => "00110", roll => "0010101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100100", store_signs_wr => '1',store_signs_addr => "010011100", load_signs_rd => '1',load_signs_addr => "010011110", min_offset => "00111", roll => "1110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100110", store_signs_wr => '1',store_signs_addr => "010011101", load_signs_rd => '1',load_signs_addr => "010011111", min_offset => "01000", roll => "0001000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101000", store_signs_wr => '1',store_signs_addr => "010011110", load_signs_rd => '1',load_signs_addr => "010100000", min_offset => "01001", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101101", store_signs_wr => '1',store_signs_addr => "010011111", load_signs_rd => '1',load_signs_addr => "010100001", min_offset => "01010", roll => "0010001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110010", store_signs_wr => '1',store_signs_addr => "010100000", load_signs_rd => '1',load_signs_addr => "010100010", min_offset => "01011", roll => "0111001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110011", store_signs_wr => '1',store_signs_addr => "010100001", load_signs_rd => '1',load_signs_addr => "010100011", min_offset => "01100", roll => "1000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000101", store_signs_wr => '1',store_signs_addr => "010100010", load_signs_rd => '1',load_signs_addr => "010100100", min_offset => "01101", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "010001", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000111", store_signs_wr => '1',store_signs_addr => "010100011", load_signs_rd => '1',load_signs_addr => "010100101", min_offset => "01110", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010111", store_signs_wr => '1',store_signs_addr => "010100100", load_signs_rd => '1',load_signs_addr => "010100110", min_offset => "00000", roll => "1111011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100101", store_signs_wr => '1',store_signs_addr => "010100101", load_signs_rd => '1',load_signs_addr => "010100111", min_offset => "00001", roll => "1111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110011", store_signs_wr => '1',store_signs_addr => "010100110", load_signs_rd => '1',load_signs_addr => "010101000", min_offset => "00010", roll => "1101011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110100", store_signs_wr => '1',store_signs_addr => "010100111", load_signs_rd => '1',load_signs_addr => "010101001", min_offset => "00011", roll => "1001110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000110", store_signs_wr => '1',store_signs_addr => "010101000", load_signs_rd => '1',load_signs_addr => "010101010", min_offset => "00100", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "010010", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000111", store_signs_wr => '1',store_signs_addr => "010101001", load_signs_rd => '1',load_signs_addr => "010101011", min_offset => "00101", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001100", store_signs_wr => '1',store_signs_addr => "010101010", load_signs_rd => '1',load_signs_addr => "010101100", min_offset => "00000", roll => "0000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001101", store_signs_wr => '1',store_signs_addr => "010101011", load_signs_rd => '1',load_signs_addr => "010101101", min_offset => "00001", roll => "1010111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001111", store_signs_wr => '1',store_signs_addr => "010101100", load_signs_rd => '1',load_signs_addr => "010101110", min_offset => "00010", roll => "0111000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010111", store_signs_wr => '1',store_signs_addr => "010101101", load_signs_rd => '1',load_signs_addr => "010101111", min_offset => "00011", roll => "1011011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110001", store_signs_wr => '1',store_signs_addr => "010101110", load_signs_rd => '1',load_signs_addr => "010110000", min_offset => "00100", roll => "0101010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110100", store_signs_wr => '1',store_signs_addr => "010101111", load_signs_rd => '1',load_signs_addr => "010110001", min_offset => "00101", roll => "0010000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110101", store_signs_wr => '1',store_signs_addr => "010110000", load_signs_rd => '1',load_signs_addr => "010110010", min_offset => "00110", roll => "0111101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000011", store_signs_wr => '1',store_signs_addr => "010110001", load_signs_rd => '1',load_signs_addr => "010110011", min_offset => "00111", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "010011", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001111", store_signs_wr => '1',store_signs_addr => "010110010", load_signs_rd => '1',load_signs_addr => "010110100", min_offset => "01000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010000", store_signs_wr => '1',store_signs_addr => "010110011", load_signs_rd => '1',load_signs_addr => "010110101", min_offset => "00000", roll => "1011100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010001", store_signs_wr => '1',store_signs_addr => "010110100", load_signs_rd => '1',load_signs_addr => "010110110", min_offset => "00001", roll => "1001100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010100", store_signs_wr => '1',store_signs_addr => "010110101", load_signs_rd => '1',load_signs_addr => "010110111", min_offset => "00010", roll => "1100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010110", store_signs_wr => '1',store_signs_addr => "010110110", load_signs_rd => '1',load_signs_addr => "010111000", min_offset => "00011", roll => "0101100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100011", store_signs_wr => '1',store_signs_addr => "010110111", load_signs_rd => '1',load_signs_addr => "010111001", min_offset => "00100", roll => "0011100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100100", store_signs_wr => '1',store_signs_addr => "010111000", load_signs_rd => '1',load_signs_addr => "010111010", min_offset => "00101", roll => "0011101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110000", store_signs_wr => '1',store_signs_addr => "010111001", load_signs_rd => '1',load_signs_addr => "010111011", min_offset => "00110", roll => "0011010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110011", store_signs_wr => '1',store_signs_addr => "010111010", load_signs_rd => '1',load_signs_addr => "010111100", min_offset => "00111", roll => "1111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110101", store_signs_wr => '1',store_signs_addr => "010111011", load_signs_rd => '1',load_signs_addr => "010111101", min_offset => "01000", roll => "0011001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110110", store_signs_wr => '1',store_signs_addr => "010111100", load_signs_rd => '1',load_signs_addr => "010111110", min_offset => "01001", roll => "0001110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000001", store_signs_wr => '1',store_signs_addr => "010111101", load_signs_rd => '1',load_signs_addr => "010111111", min_offset => "01010", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "010100", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000010", store_signs_wr => '1',store_signs_addr => "010111110", load_signs_rd => '1',load_signs_addr => "011000000", min_offset => "01011", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001001", store_signs_wr => '1',store_signs_addr => "010111111", load_signs_rd => '1',load_signs_addr => "011000001", min_offset => "00000", roll => "0010100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010010", store_signs_wr => '1',store_signs_addr => "011000000", load_signs_rd => '1',load_signs_addr => "011000010", min_offset => "00001", roll => "1011111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010110", store_signs_wr => '1',store_signs_addr => "011000001", load_signs_rd => '1',load_signs_addr => "011000011", min_offset => "00010", roll => "0010000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011100", store_signs_wr => '1',store_signs_addr => "011000010", load_signs_rd => '1',load_signs_addr => "011000100", min_offset => "00011", roll => "0111111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011110", store_signs_wr => '1',store_signs_addr => "011000011", load_signs_rd => '1',load_signs_addr => "011000101", min_offset => "00100", roll => "1101000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011111", store_signs_wr => '1',store_signs_addr => "011000100", load_signs_rd => '1',load_signs_addr => "011000110", min_offset => "00101", roll => "0010101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100100", store_signs_wr => '1',store_signs_addr => "011000101", load_signs_rd => '1',load_signs_addr => "011000111", min_offset => "00110", roll => "0101110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101101", store_signs_wr => '1',store_signs_addr => "011000110", load_signs_rd => '1',load_signs_addr => "011001000", min_offset => "00111", roll => "1001111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110011", store_signs_wr => '1',store_signs_addr => "011000111", load_signs_rd => '1',load_signs_addr => "011001001", min_offset => "01000", roll => "0001010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110110", store_signs_wr => '1',store_signs_addr => "011001000", load_signs_rd => '1',load_signs_addr => "011001010", min_offset => "01001", roll => "0111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110111", store_signs_wr => '1',store_signs_addr => "011001001", load_signs_rd => '1',load_signs_addr => "011001011", min_offset => "01010", roll => "0101011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001010", store_signs_wr => '1',store_signs_addr => "011001010", load_signs_rd => '1',load_signs_addr => "011001100", min_offset => "01011", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "010101", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001011", store_signs_wr => '1',store_signs_addr => "011001011", load_signs_rd => '1',load_signs_addr => "011001101", min_offset => "01100", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011011", store_signs_wr => '1',store_signs_addr => "011001100", load_signs_rd => '1',load_signs_addr => "011001110", min_offset => "00000", roll => "1000010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011100", store_signs_wr => '1',store_signs_addr => "011001101", load_signs_rd => '1',load_signs_addr => "011001111", min_offset => "00001", roll => "1010011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011101", store_signs_wr => '1',store_signs_addr => "011001110", load_signs_rd => '1',load_signs_addr => "011010000", min_offset => "00010", roll => "0000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011110", store_signs_wr => '1',store_signs_addr => "011001111", load_signs_rd => '1',load_signs_addr => "011010001", min_offset => "00011", roll => "1011111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100011", store_signs_wr => '1',store_signs_addr => "011010000", load_signs_rd => '1',load_signs_addr => "011010010", min_offset => "00100", roll => "1000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101010", store_signs_wr => '1',store_signs_addr => "011010001", load_signs_rd => '1',load_signs_addr => "011010011", min_offset => "00101", roll => "1100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110111", store_signs_wr => '1',store_signs_addr => "011010010", load_signs_rd => '1',load_signs_addr => "011010100", min_offset => "00110", roll => "1010100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111000", store_signs_wr => '1',store_signs_addr => "011010011", load_signs_rd => '1',load_signs_addr => "011010101", min_offset => "00111", roll => "0010101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000001", store_signs_wr => '1',store_signs_addr => "011010100", load_signs_rd => '1',load_signs_addr => "011010110", min_offset => "01000", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "010110", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000100", store_signs_wr => '1',store_signs_addr => "011010101", load_signs_rd => '1',load_signs_addr => "011010111", min_offset => "01001", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001110", store_signs_wr => '1',store_signs_addr => "011010110", load_signs_rd => '1',load_signs_addr => "011011000", min_offset => "00000", roll => "0110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010001", store_signs_wr => '1',store_signs_addr => "011010111", load_signs_rd => '1',load_signs_addr => "011011001", min_offset => "00001", roll => "1011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010010", store_signs_wr => '1',store_signs_addr => "011011000", load_signs_rd => '1',load_signs_addr => "011011010", min_offset => "00010", roll => "1110010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010111", store_signs_wr => '1',store_signs_addr => "011011001", load_signs_rd => '1',load_signs_addr => "011011011", min_offset => "00011", roll => "0011100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011011", store_signs_wr => '1',store_signs_addr => "011011010", load_signs_rd => '1',load_signs_addr => "011011100", min_offset => "00100", roll => "1001111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011111", store_signs_wr => '1',store_signs_addr => "011011011", load_signs_rd => '1',load_signs_addr => "011011101", min_offset => "00101", roll => "0001110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100011", store_signs_wr => '1',store_signs_addr => "011011100", load_signs_rd => '1',load_signs_addr => "011011110", min_offset => "00110", roll => "0100100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101101", store_signs_wr => '1',store_signs_addr => "011011101", load_signs_rd => '1',load_signs_addr => "011011111", min_offset => "00111", roll => "1011010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101111", store_signs_wr => '1',store_signs_addr => "011011110", load_signs_rd => '1',load_signs_addr => "011100000", min_offset => "01000", roll => "0010011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110011", store_signs_wr => '1',store_signs_addr => "011011111", load_signs_rd => '1',load_signs_addr => "011100001", min_offset => "01001", roll => "0101100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110101", store_signs_wr => '1',store_signs_addr => "011100000", load_signs_rd => '1',load_signs_addr => "011100010", min_offset => "01010", roll => "0110100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110111", store_signs_wr => '1',store_signs_addr => "011100001", load_signs_rd => '1',load_signs_addr => "011100011", min_offset => "01011", roll => "0011011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111000", store_signs_wr => '1',store_signs_addr => "011100010", load_signs_rd => '1',load_signs_addr => "011100100", min_offset => "01100", roll => "0101001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111001", store_signs_wr => '1',store_signs_addr => "011100011", load_signs_rd => '1',load_signs_addr => "011100101", min_offset => "01101", roll => "1100000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000010", store_signs_wr => '1',store_signs_addr => "011100100", load_signs_rd => '1',load_signs_addr => "011100110", min_offset => "01110", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "010111", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000101", store_signs_wr => '1',store_signs_addr => "011100101", load_signs_rd => '1',load_signs_addr => "011100111", min_offset => "01111", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001110", store_signs_wr => '1',store_signs_addr => "011100110", load_signs_rd => '1',load_signs_addr => "011101000", min_offset => "00000", roll => "1001000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010001", store_signs_wr => '1',store_signs_addr => "011100111", load_signs_rd => '1',load_signs_addr => "011101001", min_offset => "00001", roll => "0110110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010100", store_signs_wr => '1',store_signs_addr => "011101000", load_signs_rd => '1',load_signs_addr => "011101010", min_offset => "00010", roll => "1000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010110", store_signs_wr => '1',store_signs_addr => "011101001", load_signs_rd => '1',load_signs_addr => "011101011", min_offset => "00011", roll => "1111100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101001", store_signs_wr => '1',store_signs_addr => "011101010", load_signs_rd => '1',load_signs_addr => "011101100", min_offset => "00100", roll => "0000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101111", store_signs_wr => '1',store_signs_addr => "011101011", load_signs_rd => '1',load_signs_addr => "011101101", min_offset => "00101", roll => "0011101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110010", store_signs_wr => '1',store_signs_addr => "011101100", load_signs_rd => '1',load_signs_addr => "011101110", min_offset => "00110", roll => "1100010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110101", store_signs_wr => '1',store_signs_addr => "011101101", load_signs_rd => '1',load_signs_addr => "011101111", min_offset => "00111", roll => "1111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110110", store_signs_wr => '1',store_signs_addr => "011101110", load_signs_rd => '1',load_signs_addr => "011110000", min_offset => "01000", roll => "0011001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111000", store_signs_wr => '1',store_signs_addr => "011101111", load_signs_rd => '1',load_signs_addr => "011110001", min_offset => "01001", roll => "1101100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111001", store_signs_wr => '1',store_signs_addr => "011110000", load_signs_rd => '1',load_signs_addr => "011110010", min_offset => "01010", roll => "1010100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111010", store_signs_wr => '1',store_signs_addr => "011110001", load_signs_rd => '1',load_signs_addr => "011110011", min_offset => "01011", roll => "1111011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000010", store_signs_wr => '1',store_signs_addr => "011110010", load_signs_rd => '1',load_signs_addr => "011110100", min_offset => "01100", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "011000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000011", store_signs_wr => '1',store_signs_addr => "011110011", load_signs_rd => '1',load_signs_addr => "011110101", min_offset => "01101", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001000", store_signs_wr => '1',store_signs_addr => "011110100", load_signs_rd => '1',load_signs_addr => "011110110", min_offset => "00000", roll => "0110010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001110", store_signs_wr => '1',store_signs_addr => "011110101", load_signs_rd => '1',load_signs_addr => "011110111", min_offset => "00001", roll => "0000110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010011", store_signs_wr => '1',store_signs_addr => "011110110", load_signs_rd => '1',load_signs_addr => "011111000", min_offset => "00010", roll => "1100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010100", store_signs_wr => '1',store_signs_addr => "011110111", load_signs_rd => '1',load_signs_addr => "011111001", min_offset => "00011", roll => "0000011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010111", store_signs_wr => '1',store_signs_addr => "011111000", load_signs_rd => '1',load_signs_addr => "011111010", min_offset => "00100", roll => "0000101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011011", store_signs_wr => '1',store_signs_addr => "011111001", load_signs_rd => '1',load_signs_addr => "011111011", min_offset => "00101", roll => "0010010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100010", store_signs_wr => '1',store_signs_addr => "011111010", load_signs_rd => '1',load_signs_addr => "011111100", min_offset => "00110", roll => "0010000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100101", store_signs_wr => '1',store_signs_addr => "011111011", load_signs_rd => '1',load_signs_addr => "011111101", min_offset => "00111", roll => "1010011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110101", store_signs_wr => '1',store_signs_addr => "011111100", load_signs_rd => '1',load_signs_addr => "011111110", min_offset => "01000", roll => "1011001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110110", store_signs_wr => '1',store_signs_addr => "011111101", load_signs_rd => '1',load_signs_addr => "011111111", min_offset => "01001", roll => "0110110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110111", store_signs_wr => '1',store_signs_addr => "011111110", load_signs_rd => '1',load_signs_addr => "100000000", min_offset => "01010", roll => "0010100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111010", store_signs_wr => '1',store_signs_addr => "011111111", load_signs_rd => '1',load_signs_addr => "100000001", min_offset => "01011", roll => "1101010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111011", store_signs_wr => '1',store_signs_addr => "100000000", load_signs_rd => '1',load_signs_addr => "100000010", min_offset => "01100", roll => "0001111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000001", store_signs_wr => '1',store_signs_addr => "100000001", load_signs_rd => '1',load_signs_addr => "100000011", min_offset => "01101", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "011001", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000110", store_signs_wr => '1',store_signs_addr => "100000010", load_signs_rd => '1',load_signs_addr => "100000100", min_offset => "01110", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010011", store_signs_wr => '1',store_signs_addr => "100000011", load_signs_rd => '1',load_signs_addr => "100000101", min_offset => "00000", roll => "1101110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010100", store_signs_wr => '1',store_signs_addr => "100000100", load_signs_rd => '1',load_signs_addr => "100000110", min_offset => "00001", roll => "0111011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010101", store_signs_wr => '1',store_signs_addr => "100000101", load_signs_rd => '1',load_signs_addr => "100000111", min_offset => "00010", roll => "0101100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010110", store_signs_wr => '1',store_signs_addr => "100000110", load_signs_rd => '1',load_signs_addr => "100001000", min_offset => "00011", roll => "0010001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010111", store_signs_wr => '1',store_signs_addr => "100000111", load_signs_rd => '1',load_signs_addr => "100001001", min_offset => "00100", roll => "0011101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011011", store_signs_wr => '1',store_signs_addr => "100001000", load_signs_rd => '1',load_signs_addr => "100001010", min_offset => "00101", roll => "0101100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101000", store_signs_wr => '1',store_signs_addr => "100001001", load_signs_rd => '1',load_signs_addr => "100001011", min_offset => "00110", roll => "0110100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101001", store_signs_wr => '1',store_signs_addr => "100001010", load_signs_rd => '1',load_signs_addr => "100001100", min_offset => "00111", roll => "1010000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101101", store_signs_wr => '1',store_signs_addr => "100001011", load_signs_rd => '1',load_signs_addr => "100001101", min_offset => "01000", roll => "1000100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101111", store_signs_wr => '1',store_signs_addr => "100001100", load_signs_rd => '1',load_signs_addr => "100001110", min_offset => "01001", roll => "0010111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110101", store_signs_wr => '1',store_signs_addr => "100001101", load_signs_rd => '1',load_signs_addr => "100001111", min_offset => "01010", roll => "1010011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110110", store_signs_wr => '1',store_signs_addr => "100001110", load_signs_rd => '1',load_signs_addr => "100010000", min_offset => "01011", roll => "0011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111011", store_signs_wr => '1',store_signs_addr => "100001111", load_signs_rd => '1',load_signs_addr => "100010001", min_offset => "01100", roll => "0000100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111100", store_signs_wr => '1',store_signs_addr => "100010000", load_signs_rd => '1',load_signs_addr => "100010010", min_offset => "01101", roll => "1110001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001000", store_signs_wr => '1',store_signs_addr => "100010001", load_signs_rd => '1',load_signs_addr => "100010011", min_offset => "01110", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "011010", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001001", store_signs_wr => '1',store_signs_addr => "100010010", load_signs_rd => '1',load_signs_addr => "100010100", min_offset => "01111", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010010", store_signs_wr => '1',store_signs_addr => "100010011", load_signs_rd => '1',load_signs_addr => "100010101", min_offset => "00000", roll => "1011010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011000", store_signs_wr => '1',store_signs_addr => "100010100", load_signs_rd => '1',load_signs_addr => "100010110", min_offset => "00001", roll => "0000011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011001", store_signs_wr => '1',store_signs_addr => "100010101", load_signs_rd => '1',load_signs_addr => "100010111", min_offset => "00010", roll => "1011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100100", store_signs_wr => '1',store_signs_addr => "100010110", load_signs_rd => '1',load_signs_addr => "100011000", min_offset => "00011", roll => "0111101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101111", store_signs_wr => '1',store_signs_addr => "100010111", load_signs_rd => '1',load_signs_addr => "100011001", min_offset => "00100", roll => "1011011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110110", store_signs_wr => '1',store_signs_addr => "100011000", load_signs_rd => '1',load_signs_addr => "100011010", min_offset => "00101", roll => "0110100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111100", store_signs_wr => '1',store_signs_addr => "100011001", load_signs_rd => '1',load_signs_addr => "100011011", min_offset => "00110", roll => "1100010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111101", store_signs_wr => '1',store_signs_addr => "100011010", load_signs_rd => '1',load_signs_addr => "100011100", min_offset => "00111", roll => "1011001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001100", store_signs_wr => '1',store_signs_addr => "100011011", load_signs_rd => '1',load_signs_addr => "100011101", min_offset => "01000", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "011011", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010111", store_signs_wr => '1',store_signs_addr => "100011100", load_signs_rd => '1',load_signs_addr => "100011110", min_offset => "01001", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011000", store_signs_wr => '1',store_signs_addr => "100011101", load_signs_rd => '1',load_signs_addr => "100011111", min_offset => "00000", roll => "0110111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011100", store_signs_wr => '1',store_signs_addr => "100011110", load_signs_rd => '1',load_signs_addr => "100100000", min_offset => "00001", roll => "0000110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100000", store_signs_wr => '1',store_signs_addr => "100011111", load_signs_rd => '1',load_signs_addr => "100100001", min_offset => "00010", roll => "1100111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101000", store_signs_wr => '1',store_signs_addr => "100100000", load_signs_rd => '1',load_signs_addr => "100100010", min_offset => "00011", roll => "0010110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101100", store_signs_wr => '1',store_signs_addr => "100100001", load_signs_rd => '1',load_signs_addr => "100100011", min_offset => "00100", roll => "0100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101110", store_signs_wr => '1',store_signs_addr => "100100010", load_signs_rd => '1',load_signs_addr => "100100100", min_offset => "00101", roll => "0011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101111", store_signs_wr => '1',store_signs_addr => "100100011", load_signs_rd => '1',load_signs_addr => "100100101", min_offset => "00110", roll => "1101000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111001", store_signs_wr => '1',store_signs_addr => "100100100", load_signs_rd => '1',load_signs_addr => "100100110", min_offset => "00111", roll => "1100000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111101", store_signs_wr => '1',store_signs_addr => "100100101", load_signs_rd => '1',load_signs_addr => "100100111", min_offset => "01000", roll => "1001000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111110", store_signs_wr => '1',store_signs_addr => "100100110", load_signs_rd => '1',load_signs_addr => "100101000", min_offset => "01001", roll => "1001011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000001", store_signs_wr => '1',store_signs_addr => "100100111", load_signs_rd => '1',load_signs_addr => "100101001", min_offset => "01010", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "011100", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001011", store_signs_wr => '1',store_signs_addr => "100101000", load_signs_rd => '1',load_signs_addr => "100101010", min_offset => "01011", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001101", store_signs_wr => '1',store_signs_addr => "100101001", load_signs_rd => '1',load_signs_addr => "100101011", min_offset => "00000", roll => "1000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010000", store_signs_wr => '1',store_signs_addr => "100101010", load_signs_rd => '1',load_signs_addr => "100101100", min_offset => "00001", roll => "1110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010010", store_signs_wr => '1',store_signs_addr => "100101011", load_signs_rd => '1',load_signs_addr => "100101101", min_offset => "00010", roll => "1010100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010110", store_signs_wr => '1',store_signs_addr => "100101100", load_signs_rd => '1',load_signs_addr => "100101110", min_offset => "00011", roll => "0000011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011000", store_signs_wr => '1',store_signs_addr => "100101101", load_signs_rd => '1',load_signs_addr => "100101111", min_offset => "00100", roll => "1010010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100011", store_signs_wr => '1',store_signs_addr => "100101110", load_signs_rd => '1',load_signs_addr => "100110000", min_offset => "00101", roll => "1011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101001", store_signs_wr => '1',store_signs_addr => "100101111", load_signs_rd => '1',load_signs_addr => "100110001", min_offset => "00110", roll => "0111100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101010", store_signs_wr => '1',store_signs_addr => "100110000", load_signs_rd => '1',load_signs_addr => "100110010", min_offset => "00111", roll => "0111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101101", store_signs_wr => '1',store_signs_addr => "100110001", load_signs_rd => '1',load_signs_addr => "100110011", min_offset => "01000", roll => "0110000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111100", store_signs_wr => '1',store_signs_addr => "100110010", load_signs_rd => '1',load_signs_addr => "100110100", min_offset => "01001", roll => "0110100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111110", store_signs_wr => '1',store_signs_addr => "100110011", load_signs_rd => '1',load_signs_addr => "100110101", min_offset => "01010", roll => "1000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111111", store_signs_wr => '1',store_signs_addr => "100110100", load_signs_rd => '1',load_signs_addr => "100110110", min_offset => "01011", roll => "1100010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000100", store_signs_wr => '1',store_signs_addr => "100110101", load_signs_rd => '1',load_signs_addr => "100110111", min_offset => "01100", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "011101", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000111", store_signs_wr => '1',store_signs_addr => "100110110", load_signs_rd => '1',load_signs_addr => "100111000", min_offset => "01101", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001010", store_signs_wr => '1',store_signs_addr => "100110111", load_signs_rd => '1',load_signs_addr => "100111001", min_offset => "00000", roll => "1000010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001111", store_signs_wr => '1',store_signs_addr => "100111000", load_signs_rd => '1',load_signs_addr => "100111010", min_offset => "00001", roll => "1100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0010000", store_signs_wr => '1',store_signs_addr => "100111001", load_signs_rd => '1',load_signs_addr => "100111011", min_offset => "00010", roll => "1110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0011101", store_signs_wr => '1',store_signs_addr => "100111010", load_signs_rd => '1',load_signs_addr => "100111100", min_offset => "00011", roll => "0001001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100001", store_signs_wr => '1',store_signs_addr => "100111011", load_signs_rd => '1',load_signs_addr => "100111101", min_offset => "00100", roll => "0111001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101000", store_signs_wr => '1',store_signs_addr => "100111100", load_signs_rd => '1',load_signs_addr => "100111110", min_offset => "00101", roll => "1000011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110000", store_signs_wr => '1',store_signs_addr => "100111101", load_signs_rd => '1',load_signs_addr => "100111111", min_offset => "00110", roll => "0000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110010", store_signs_wr => '1',store_signs_addr => "100111110", load_signs_rd => '1',load_signs_addr => "101000000", min_offset => "00111", roll => "0010011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111111", store_signs_wr => '1',store_signs_addr => "100111111", load_signs_rd => '1',load_signs_addr => "101000001", min_offset => "01000", roll => "0001000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "1000000", store_signs_wr => '1',store_signs_addr => "101000000", load_signs_rd => '1',load_signs_addr => "101000010", min_offset => "01001", roll => "1111001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000010", store_signs_wr => '1',store_signs_addr => "101000001", load_signs_rd => '1',load_signs_addr => "101000011", min_offset => "01010", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "011110", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000100", store_signs_wr => '1',store_signs_addr => "101000010", load_signs_rd => '1',load_signs_addr => "101000100", min_offset => "01011", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000110", store_signs_wr => '1',store_signs_addr => "101000011", load_signs_rd => '1',load_signs_addr => "101000101", min_offset => "00000", roll => "0110000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001000", store_signs_wr => '1',store_signs_addr => "101000100", load_signs_rd => '1',load_signs_addr => "101000110", min_offset => "00001", roll => "0010110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100001", store_signs_wr => '1',store_signs_addr => "101000101", load_signs_rd => '1',load_signs_addr => "101000111", min_offset => "00010", roll => "0100100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101001", store_signs_wr => '1',store_signs_addr => "101000110", load_signs_rd => '1',load_signs_addr => "101001000", min_offset => "00011", roll => "0110001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101010", store_signs_wr => '1',store_signs_addr => "101000111", load_signs_rd => '1',load_signs_addr => "101001001", min_offset => "00100", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101011", store_signs_wr => '1',store_signs_addr => "101001000", load_signs_rd => '1',load_signs_addr => "101001010", min_offset => "00101", roll => "0011010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101111", store_signs_wr => '1',store_signs_addr => "101001001", load_signs_rd => '1',load_signs_addr => "101001011", min_offset => "00110", roll => "0000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110010", store_signs_wr => '1',store_signs_addr => "101001010", load_signs_rd => '1',load_signs_addr => "101001100", min_offset => "00111", roll => "0110000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110100", store_signs_wr => '1',store_signs_addr => "101001011", load_signs_rd => '1',load_signs_addr => "101001101", min_offset => "01000", roll => "0010110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111000", store_signs_wr => '1',store_signs_addr => "101001100", load_signs_rd => '1',load_signs_addr => "101001110", min_offset => "01001", roll => "0011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111001", store_signs_wr => '1',store_signs_addr => "101001101", load_signs_rd => '1',load_signs_addr => "101001111", min_offset => "01010", roll => "0100001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111010", store_signs_wr => '1',store_signs_addr => "101001110", load_signs_rd => '1',load_signs_addr => "101010000", min_offset => "01011", roll => "1100111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111100", store_signs_wr => '1',store_signs_addr => "101001111", load_signs_rd => '1',load_signs_addr => "101010001", min_offset => "01100", roll => "1100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111101", store_signs_wr => '1',store_signs_addr => "101010000", load_signs_rd => '1',load_signs_addr => "101010010", min_offset => "01101", roll => "1100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "1000000", store_signs_wr => '1',store_signs_addr => "101010001", load_signs_rd => '1',load_signs_addr => "101010011", min_offset => "01110", roll => "1000101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "1000001", store_signs_wr => '1',store_signs_addr => "101010010", load_signs_rd => '1',load_signs_addr => "101010100", min_offset => "01111", roll => "1000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0000011", store_signs_wr => '1',store_signs_addr => "101010011", load_signs_rd => '1',load_signs_addr => "101010101", min_offset => "10000", roll => "0000000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "011111", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001000", store_signs_wr => '1',store_signs_addr => "101010100", load_signs_rd => '1',load_signs_addr => "101010110", min_offset => "10001", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0001101", store_signs_wr => '1',store_signs_addr => "101010101", load_signs_rd => '1',load_signs_addr => "101010111", min_offset => "00000", roll => "1111100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0100001", store_signs_wr => '1',store_signs_addr => "101010110", load_signs_rd => '1',load_signs_addr => "101011000", min_offset => "00001", roll => "1000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101010", store_signs_wr => '1',store_signs_addr => "101010111", load_signs_rd => '1',load_signs_addr => "101011001", min_offset => "00010", roll => "1011111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101100", store_signs_wr => '1',store_signs_addr => "101011000", load_signs_rd => '1',load_signs_addr => "101011010", min_offset => "00011", roll => "0000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0101110", store_signs_wr => '1',store_signs_addr => "101011001", load_signs_rd => '1',load_signs_addr => "101011011", min_offset => "00100", roll => "0100111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0110110", store_signs_wr => '1',store_signs_addr => "101011010", load_signs_rd => '1',load_signs_addr => "101011100", min_offset => "00101", roll => "1110100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "0111011", store_signs_wr => '1',store_signs_addr => "101011011", load_signs_rd => '1',load_signs_addr => "101011101", min_offset => "00110", roll => "1000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '1',load_vn_addr => "1000001", store_signs_wr => '1',store_signs_addr => "101011100", load_signs_rd => '1',load_signs_addr => "101011110", min_offset => "00111", roll => "0010000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '1',store_signs_addr => "101011101", load_signs_rd => '1',load_signs_addr => "000000000", min_offset => "01000", roll => "1101010")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "0000001", result_wr => '0',result_addr => "0000000", store_cn_wr => '1',store_cn_addr => "100000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '1',store_signs_addr => "101011110", load_signs_rd => '1',load_signs_addr => "001010100", min_offset => "01001", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000000001", min_offset => "00000", roll => "1100101")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '1',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000100011", min_offset => "00000", roll => "0101010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001010101", min_offset => "00000", roll => "1001101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010111111", min_offset => "00000", roll => "1001100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011010110", min_offset => "00000", roll => "1000010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100000011", min_offset => "00000", roll => "0010100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0000010", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100101001", min_offset => "00000", roll => "0110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0000001", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000111101", min_offset => "00000", roll => "1101110")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '1',store_vn_addr => "0000001", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001001000", min_offset => "00000", roll => "1000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001010110", min_offset => "00000", roll => "1000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001101111", min_offset => "00000", roll => "0110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010000001", min_offset => "00000", roll => "1101111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011000000", min_offset => "00000", roll => "1011001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011100110", min_offset => "00000", roll => "1000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011110100", min_offset => "00000", roll => "1011111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0000011", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101000011", min_offset => "00000", roll => "1001000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0000010", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000100100", min_offset => "00000", roll => "0110010")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '1',store_vn_addr => "0000010", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010010101", min_offset => "00000", roll => "0110000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010110011", min_offset => "00000", roll => "0001110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011110101", min_offset => "00000", roll => "0111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0000100", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101010101", min_offset => "00000", roll => "1011100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0000011", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001110111", min_offset => "00000", roll => "0000110")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '1',store_vn_addr => "0000011", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010010110", min_offset => "00000", roll => "1111100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011010111", min_offset => "00000", roll => "1100000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100110111", min_offset => "00000", roll => "1110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0000101", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101000100", min_offset => "00000", roll => "1011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0000100", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000100101", min_offset => "00000", roll => "1000010")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '1',store_vn_addr => "0000100", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000110000", min_offset => "00000", roll => "0010110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010000010", min_offset => "00000", roll => "0110001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010100100", min_offset => "00000", roll => "0011111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0000110", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011100111", min_offset => "00000", roll => "0001001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0000101", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001110000", min_offset => "00000", roll => "1111011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '1',store_vn_addr => "0000101", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010101010", min_offset => "00000", roll => "0110110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100000100", min_offset => "00000", roll => "1000101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0000111", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101000101", min_offset => "00000", roll => "0000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0000110", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000011000", min_offset => "00000", roll => "0111011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '1',store_vn_addr => "0000110", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000110001", min_offset => "00000", roll => "0100100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001011101", min_offset => "00000", roll => "1110000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001110001", min_offset => "00000", roll => "0110010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001111000", min_offset => "00000", roll => "0000010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010010111", min_offset => "00000", roll => "1011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010100101", min_offset => "00000", roll => "0111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010101011", min_offset => "00000", roll => "0110110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0001000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100111000", min_offset => "00000", roll => "1111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0000111", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000000101", min_offset => "00000", roll => "1010111")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '1',store_vn_addr => "0000111", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000001100", min_offset => "00000", roll => "1100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000011001", min_offset => "00000", roll => "0010110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010011000", min_offset => "00000", roll => "1010111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011110110", min_offset => "00000", roll => "1001111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100010011", min_offset => "00000", roll => "0100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101000110", min_offset => "00000", roll => "1100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0001001", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101010110", min_offset => "00000", roll => "1011010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0001000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000100110", min_offset => "00000", roll => "0110001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '1',store_vn_addr => "0001000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010000011", min_offset => "00000", roll => "1000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011000001", min_offset => "00000", roll => "1111000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0001010", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100010100", min_offset => "00000", roll => "1000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0001001", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000000110", min_offset => "00000", roll => "0010000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '1',store_vn_addr => "0001001", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001001001", min_offset => "00000", roll => "0000011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001111001", min_offset => "00000", roll => "1011010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011001100", min_offset => "00000", roll => "0111100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0001011", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100111001", min_offset => "00000", roll => "0000110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0001010", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000100111", min_offset => "00000", roll => "1000010")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '1',store_vn_addr => "0001010", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000111110", min_offset => "00000", roll => "1110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011001101", min_offset => "00000", roll => "1110110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0001100", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100101010", min_offset => "00000", roll => "0101001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0001011", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000000111", min_offset => "00000", roll => "1010011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '1',store_vn_addr => "0001011", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000110010", min_offset => "00000", roll => "1110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001010111", min_offset => "00000", roll => "1011110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010000100", min_offset => "00000", roll => "0001111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010101100", min_offset => "00000", roll => "0110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0001101", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100011101", min_offset => "00000", roll => "1011011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0001100", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000001000", min_offset => "00000", roll => "0111000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '1',store_vn_addr => "0001100", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000001101", min_offset => "00000", roll => "0110111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000101000", min_offset => "00000", roll => "0001000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000110011", min_offset => "00000", roll => "0110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001011110", min_offset => "00000", roll => "1110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001111010", min_offset => "00000", roll => "0111111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010101101", min_offset => "00000", roll => "1101001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100101011", min_offset => "00000", roll => "1101111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0001110", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101010111", min_offset => "00000", roll => "1011011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0001101", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000111111", min_offset => "00000", roll => "1010100")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '1',store_vn_addr => "0001101", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001001010", min_offset => "00000", roll => "1011111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001100111", min_offset => "00000", roll => "1001100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010000101", min_offset => "00000", roll => "0101110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010001111", min_offset => "00000", roll => "0110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011011000", min_offset => "00000", roll => "0111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011101000", min_offset => "00000", roll => "1110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0001111", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011110111", min_offset => "00000", roll => "1110010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0001110", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000010010", min_offset => "00000", roll => "1000111")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '1',store_vn_addr => "0001110", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000011101", min_offset => "00000", roll => "0000011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001000000", min_offset => "00000", roll => "1000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001110010", min_offset => "00000", roll => "0111111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010101110", min_offset => "00000", roll => "0101111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010110100", min_offset => "00000", roll => "1011111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0010000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100111010", min_offset => "00000", roll => "0101010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0001111", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000110100", min_offset => "00000", roll => "1001100")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '1',store_vn_addr => "0001111", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001111011", min_offset => "00000", roll => "0001001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010110101", min_offset => "00000", roll => "0000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100101100", min_offset => "00000", roll => "0110011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0010001", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100111011", min_offset => "00000", roll => "1100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0010000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001001011", min_offset => "00000", roll => "0000011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '1',store_vn_addr => "0010000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010110110", min_offset => "00000", roll => "0111001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011011001", min_offset => "00000", roll => "1001011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0010010", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011101001", min_offset => "00000", roll => "0101100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0010001", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000110101", min_offset => "00000", roll => "0011100")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '1',store_vn_addr => "0010001", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001001100", min_offset => "00000", roll => "1111100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001111100", min_offset => "00000", roll => "0000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010000110", min_offset => "00000", roll => "0100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011000010", min_offset => "00000", roll => "0100111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011011010", min_offset => "00000", roll => "0010010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100010101", min_offset => "00000", roll => "0111111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0010011", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100101101", min_offset => "00000", roll => "1001111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0010010", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000010011", min_offset => "00000", roll => "1011000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000100", store_vn_wr => '1',store_vn_addr => "0010010", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000011010", min_offset => "00000", roll => "1010010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000101001", min_offset => "00000", roll => "1000101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001000001", min_offset => "00000", roll => "1000011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011111000", min_offset => "00000", roll => "1100010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0010100", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100000101", min_offset => "00000", roll => "1101101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0010011", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001101000", min_offset => "00000", roll => "0000101")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '1',store_vn_addr => "0010011", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001111101", min_offset => "00000", roll => "0101100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010011001", min_offset => "00000", roll => "1000011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010110111", min_offset => "00000", roll => "0111001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011101010", min_offset => "00000", roll => "0100111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011111001", min_offset => "00000", roll => "0011100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0010101", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100000110", min_offset => "00000", roll => "0000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0010110", result_wr => '1',result_addr => "0010100", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100000111", min_offset => "00000", roll => "0010010")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0010101", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '1',store_vn_addr => "0010100", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000011110", min_offset => "00000", roll => "0010001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '1',store_vn_addr => "0010101", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000110110", min_offset => "00000", roll => "0011101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010011010", min_offset => "00000", roll => "0111011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010111000", min_offset => "00000", roll => "1100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011000011", min_offset => "00000", roll => "1011100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011101011", min_offset => "00000", roll => "0011101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100001000", min_offset => "00000", roll => "1101000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0010111", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100101110", min_offset => "00000", roll => "0011101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0010110", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000110111", min_offset => "00000", roll => "0101100")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '1',store_vn_addr => "0010110", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010000111", min_offset => "00000", roll => "1011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010100110", min_offset => "00000", roll => "1100011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010101111", min_offset => "00000", roll => "0100111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011011011", min_offset => "00000", roll => "1101011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011111010", min_offset => "00000", roll => "0010000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100001001", min_offset => "00000", roll => "0001110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0011000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100011110", min_offset => "00000", roll => "0010000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0010111", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010001000", min_offset => "00000", roll => "0110100")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '1',store_vn_addr => "0010111", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100010110", min_offset => "00000", roll => "0000110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100011111", min_offset => "00000", roll => "1000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0011001", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100101111", min_offset => "00000", roll => "0111101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0011000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000101010", min_offset => "00000", roll => "1100111")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '1',store_vn_addr => "0011000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001000010", min_offset => "00000", roll => "0111100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001001101", min_offset => "00000", roll => "1111001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001011111", min_offset => "00000", roll => "0111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010001001", min_offset => "00000", roll => "0111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0011010", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100010111", min_offset => "00000", roll => "1111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0011001", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000000010", min_offset => "00000", roll => "0000100")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '1',store_vn_addr => "0011001", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000001001", min_offset => "00000", roll => "1011011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000011111", min_offset => "00000", roll => "1111011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001000011", min_offset => "00000", roll => "0111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0011011", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001100000", min_offset => "00000", roll => "0101111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0011010", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000001110", min_offset => "00000", roll => "1110000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '1',store_vn_addr => "0011010", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000010100", min_offset => "00000", roll => "1001001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000100000", min_offset => "00000", roll => "1010111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001000100", min_offset => "00000", roll => "1111000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001001110", min_offset => "00000", roll => "1000101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001101001", min_offset => "00000", roll => "1110100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010011011", min_offset => "00000", roll => "1010011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011001110", min_offset => "00000", roll => "1000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011011100", min_offset => "00000", roll => "0010101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011111011", min_offset => "00000", roll => "0000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0011100", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100001010", min_offset => "00000", roll => "0100100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0011011", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000000011", min_offset => "00000", roll => "1010011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '1',store_vn_addr => "0011011", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011000100", min_offset => "00000", roll => "1010000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011001111", min_offset => "00000", roll => "1011100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0011101", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100100000", min_offset => "00000", roll => "0010101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0011100", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000001111", min_offset => "00000", roll => "1011111")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '1',store_vn_addr => "0011100", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000101011", min_offset => "00000", roll => "0010110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001000101", min_offset => "00000", roll => "1110010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010011100", min_offset => "00000", roll => "1001011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011010000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0011110", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100111100", min_offset => "00000", roll => "1110101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0011101", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001011000", min_offset => "00000", roll => "1000001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '1',store_vn_addr => "0011101", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001100001", min_offset => "00000", roll => "1000011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010010000", min_offset => "00000", roll => "0101001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010011101", min_offset => "00000", roll => "1000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011000101", min_offset => "00000", roll => "1000010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0011111", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011010001", min_offset => "00000", roll => "0001000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0011110", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001001111", min_offset => "00000", roll => "0101110")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '1',store_vn_addr => "0011110", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001011001", min_offset => "00000", roll => "1100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001100010", min_offset => "00000", roll => "1101101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011000110", min_offset => "00000", roll => "1110000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0100000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011011101", min_offset => "00000", roll => "1010111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0011111", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000010101", min_offset => "00000", roll => "1001111")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '1',store_vn_addr => "0011111", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000101100", min_offset => "00000", roll => "1011010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000111000", min_offset => "00000", roll => "1101011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001100011", min_offset => "00000", roll => "1101011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001110011", min_offset => "00000", roll => "1100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010001010", min_offset => "00000", roll => "1100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0100001", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100100001", min_offset => "00000", roll => "0101101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0100000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100111101", min_offset => "00000", roll => "0010100")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '1',store_vn_addr => "0100000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101000111", min_offset => "00000", roll => "0100110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0100010", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101011000", min_offset => "00000", roll => "0000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0100001", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000000100", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '1',store_vn_addr => "0100001", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000001010", min_offset => "00000", roll => "0000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000111001", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010001011", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0100011", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011111100", min_offset => "00000", roll => "1110001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0100010", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000001011", min_offset => "00000", roll => "1011110")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '1',store_vn_addr => "0100010", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000010000", min_offset => "00000", roll => "1011001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001111110", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010111001", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011010010", min_offset => "00000", roll => "0010110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011011110", min_offset => "00000", roll => "0011010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0100100", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100110000", min_offset => "00000", roll => "1010100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0100011", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000010001", min_offset => "00000", roll => "0010011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '1',store_vn_addr => "0100011", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000010110", min_offset => "00000", roll => "0111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001100100", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010011110", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010111010", min_offset => "00000", roll => "0100001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011000111", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0100101", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100011000", min_offset => "00000", roll => "1111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0100100", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000010111", min_offset => "00000", roll => "0001010")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000100", store_vn_wr => '1',store_vn_addr => "0100100", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000011011", min_offset => "00000", roll => "0110100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001010000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001101010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010001100", min_offset => "00000", roll => "0110001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010100111", min_offset => "00000", roll => "1110110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0100110", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011111101", min_offset => "00000", roll => "1010011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0100101", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000011100", min_offset => "00000", roll => "1001110")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '1',store_vn_addr => "0100101", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000100001", min_offset => "00000", roll => "0110110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000101101", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000111010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001101011", min_offset => "00000", roll => "0000010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0100111", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010011111", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0100110", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000100010", min_offset => "00000", roll => "1111101")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '1',store_vn_addr => "0100110", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000101110", min_offset => "00000", roll => "0010001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001011010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0101000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010010001", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0100111", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000101111", min_offset => "00000", roll => "0101100")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '1',store_vn_addr => "0100111", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000111011", min_offset => "00000", roll => "0100100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010100000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100001011", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100100010", min_offset => "00000", roll => "0111001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0101001", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100111110", min_offset => "00000", roll => "1000100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0101000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "000111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "000111100", min_offset => "00000", roll => "0011000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '1',store_vn_addr => "0101000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001000110", min_offset => "00000", roll => "0010011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001010001", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001110100", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011101100", min_offset => "00000", roll => "0110111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100001100", min_offset => "00000", roll => "0111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100110001", min_offset => "00000", roll => "1100010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0101010", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101001000", min_offset => "00000", roll => "0010111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0101001", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001000111", min_offset => "00000", roll => "0110000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '1',store_vn_addr => "0101001", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001010010", min_offset => "00000", roll => "0011010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011010011", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100110010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101001001", min_offset => "00000", roll => "0010101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0101011", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101011001", min_offset => "00000", roll => "0110100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0101010", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001010011", min_offset => "00000", roll => "0000001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '1',store_vn_addr => "0101010", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001011011", min_offset => "00000", roll => "0100111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0101100", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101001010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0101011", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001011100", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '1',store_vn_addr => "0101011", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001100101", min_offset => "00000", roll => "0110000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001101100", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100100011", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0101101", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101011010", min_offset => "00000", roll => "1001101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0101100", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001100110", min_offset => "00000", roll => "1101000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '1',store_vn_addr => "0101100", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001101101", min_offset => "00000", roll => "1110100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010100001", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011001000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011011111", min_offset => "00000", roll => "1000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100001101", min_offset => "00000", roll => "0111110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0101110", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100110011", min_offset => "00000", roll => "0101100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0101101", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001101110", min_offset => "00000", roll => "1010011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '1',store_vn_addr => "0101101", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001110101", min_offset => "00000", roll => "1000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100100100", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0101111", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101011011", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0101110", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001110110", min_offset => "00000", roll => "1100000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '1',store_vn_addr => "0101110", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "001111111", min_offset => "00000", roll => "1000111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011100000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011101101", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100001110", min_offset => "00000", roll => "0110100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100011001", min_offset => "00000", roll => "1111010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100100101", min_offset => "00000", roll => "0011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0110000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101001011", min_offset => "00000", roll => "1100010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0101111", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010000000", min_offset => "00000", roll => "1001000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '1',store_vn_addr => "0101111", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010001101", min_offset => "00000", roll => "0010110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010010010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010111011", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0110001", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100111111", min_offset => "00000", roll => "0101011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0110000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "001111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010001110", min_offset => "00000", roll => "0011001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '1',store_vn_addr => "0110000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010010011", min_offset => "00000", roll => "0001000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0110010", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010110000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0110001", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010010100", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '1',store_vn_addr => "0110001", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010100010", min_offset => "00000", roll => "0111101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011101110", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101000000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0110011", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101001100", min_offset => "00000", roll => "0011001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0110010", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010100011", min_offset => "00000", roll => "1111001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '1',store_vn_addr => "0110010", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010101000", min_offset => "00000", roll => "0011000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010111100", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011001001", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0110100", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011100001", min_offset => "00000", roll => "0001110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0110011", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010101001", min_offset => "00000", roll => "0101011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '1',store_vn_addr => "0110011", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010110001", min_offset => "00000", roll => "0011011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0110101", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101001101", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0110100", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010110010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '1',store_vn_addr => "0110100", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010111101", min_offset => "00000", roll => "0100001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011100010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011101111", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011111110", min_offset => "00000", roll => "0101001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0110110", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100001111", min_offset => "00000", roll => "1101100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0110101", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "010111110", min_offset => "00000", roll => "0010100")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '1',store_vn_addr => "0110101", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011001010", min_offset => "00000", roll => "0000100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011110000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011111111", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100010000", min_offset => "00000", roll => "1010100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100011010", min_offset => "00000", roll => "1101010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0110111", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101011100", min_offset => "00000", roll => "1110001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0110110", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011001011", min_offset => "00000", roll => "1011001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '1',store_vn_addr => "0110110", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011010100", min_offset => "00000", roll => "0010000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011100011", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0111000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100000000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0110111", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011010101", min_offset => "00000", roll => "1100000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '1',store_vn_addr => "0110111", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011100100", min_offset => "00000", roll => "0001111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011110001", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0111001", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101001110", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0111000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "010111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011100101", min_offset => "00000", roll => "1111011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '1',store_vn_addr => "0111000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011110010", min_offset => "00000", roll => "1100111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100100110", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0111010", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101001111", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0111001", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "011110011", min_offset => "00000", roll => "1001011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '1',store_vn_addr => "0111001", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100000001", min_offset => "00000", roll => "1100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0111011", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101010000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0111010", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011001", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100000010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '1',store_vn_addr => "0111010", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100010001", min_offset => "00000", roll => "1100101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0111100", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101011101", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0111011", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011010", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100010010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '1',store_vn_addr => "0111011", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100011011", min_offset => "00000", roll => "1101010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100110100", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0111101", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101010001", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0111100", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011011", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100011100", min_offset => "00000", roll => "1100010")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '1',store_vn_addr => "0111100", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100100111", min_offset => "00000", roll => "1000101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "0111110", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101010010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0111101", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011100", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100101000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "0111111", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '1',store_vn_addr => "0111101", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100110101", min_offset => "00000", roll => "1000001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0111110", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011101", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "100110110", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "1000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '1',store_vn_addr => "0111110", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101000001", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "0111111", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011110", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101000010", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "1000001", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '1',store_vn_addr => "0111111", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101010011", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "1000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "011111", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101010100", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '1',load_cn_addr => "100000", store_vn_wr => '1',store_vn_addr => "1000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '1',load_signs_addr => "101011110", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '1',result_addr => "1000001", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '0',load_cn_addr => "000000", store_vn_wr => '0',store_vn_addr => "0000000", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '0',load_signs_addr => "000000000", min_offset => "00000", roll => "0000000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "0000000", result_wr => '0',result_addr => "0000000", store_cn_wr => '0',store_cn_addr => "000000", load_cn_rd => '0',load_cn_addr => "000000", store_vn_wr => '1',store_vn_addr => "1000001", load_vn_rd => '0',load_vn_addr => "0000000", store_signs_wr => '0',store_signs_addr => "000000000", load_signs_rd => '0',load_signs_addr => "000000000", min_offset => "00000", roll => "0000000")));
end package;
package body common is
function pack(int_in : inst_t) return std_logic_vector is
variable rv : vec_inst_t;
begin
rv(1-1) := int_in.row_end;
rv(2-1) := int_in.col_end;
rv(3-1) := int_in.llr_mem_rd;
rv(10-1 downto 3) := std_logic_vector(int_in.llr_mem_addr);
rv(17-1 downto 10) := std_logic_vector(int_in.result_addr);
rv(18-1) := int_in.result_wr;
rv(19-1) := int_in.store_cn_wr;
rv(25-1 downto 19) := std_logic_vector(int_in.store_cn_addr);
rv(26-1) := int_in.load_cn_rd;
rv(32-1 downto 26) := std_logic_vector(int_in.load_cn_addr);
rv(33-1) := int_in.store_vn_wr;
rv(40-1 downto 33) := std_logic_vector(int_in.store_vn_addr);
rv(41-1) := int_in.load_vn_rd;
rv(48-1 downto 41) := std_logic_vector(int_in.load_vn_addr);
rv(49-1) := int_in.store_signs_wr;
rv(58-1 downto 49) := std_logic_vector(int_in.store_signs_addr);
rv(59-1) := int_in.load_signs_rd;
rv(68-1 downto 59) := std_logic_vector(int_in.load_signs_addr);
rv(73-1 downto 68) := std_logic_vector(int_in.min_offset);
rv(80-1 downto 73) := std_logic_vector(int_in.roll);
return rv;
end function;
function unpack(int_in : std_logic_vector) return inst_t is
variable rv : inst_t;
begin
rv.row_end:= (int_in(1-1));
rv.col_end:= (int_in(2-1));
rv.llr_mem_rd:= (int_in(3-1));
rv.llr_mem_addr:= unsigned(int_in(10-1 downto 3));
rv.result_addr:= unsigned(int_in(17-1 downto 10));
rv.result_wr:= (int_in(18-1));
rv.store_cn_wr:= (int_in(19-1));
rv.store_cn_addr:= unsigned(int_in(25-1 downto 19));
rv.load_cn_rd:= (int_in(26-1));
rv.load_cn_addr:= unsigned(int_in(32-1 downto 26));
rv.store_vn_wr:= (int_in(33-1));
rv.store_vn_addr:= unsigned(int_in(40-1 downto 33));
rv.load_vn_rd:= (int_in(41-1));
rv.load_vn_addr:= unsigned(int_in(48-1 downto 41));
rv.store_signs_wr:= (int_in(49-1));
rv.store_signs_addr:= unsigned(int_in(58-1 downto 49));
rv.load_signs_rd:= (int_in(59-1));
rv.load_signs_addr:= unsigned(int_in(68-1 downto 59));
rv.min_offset:= unsigned(int_in(73-1 downto 68));
rv.roll:= unsigned(int_in(80-1 downto 73));
return rv;
end function;
end package body;
