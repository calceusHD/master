
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;

package common is
constant RNG_WORDS : natural := 11;
constant ENCODE_BITS_IN : natural := 324;
constant ENCODE_BITS_OUT : natural := 648;
constant ENCODE_SLAVE_PADDING : natural := 352;
constant ENCODE_MASTER_PADDING : natural := 8;
constant BIT_SLAVE_PADDING : natural := 26;
constant BIT_MASTER_PADDING : natural := 24;
constant DECODE_SLAVE_PADDING : natural := 8;
constant DECODE_MASTER_PADDING : natural := 8;
constant LLR_BITS : natural := 7;
type llr_row_t is array(0 to 1-1) of signed(7-1 downto 0);
type llr_array_t is array(0 to 27-1, 0  to 1-1) of signed(7-1 downto 0);
type llr_column_t is array(0 to 27-1) of signed(7-1 downto 0);
subtype column_sum_t is signed(11-1 downto 0);
type column_sum_array_t is array(0 to 27-1) of column_sum_t;
subtype min_signs_t is std_logic_vector(0 to 27-1);
subtype min_t is unsigned(7-1 downto 0);
type min_array_t is array(0 to 27-1) of unsigned(7-1 downto 0);
type signs_t is array(0 to 27-1) of std_logic_vector(0 to 1-1);
subtype min_id_t is unsigned(3-1 downto 0);
type min_id_array_t is array(0 to 27-1) of min_id_t;
type roll_count_t is array(0 to 1-1) of natural;
subtype row_addr_t is unsigned(5-1 downto 0);
subtype col_addr_t is unsigned(4-1 downto 0);
subtype signs_addr_t is unsigned(7-1 downto 0);
subtype roll_t is unsigned(5-1 downto 0);
constant ROLL_COUNT : roll_count_t := (0, others => 0);
constant HQC_COLUMNS : natural := 24;
constant VN_MEM_BITS : natural := 5;
constant CN_MEM_BITS : natural := 4;
subtype vec_inst_t is std_logic_vector(60-1 downto 0);
type inst_t is 
    record
        row_end : std_logic;
        col_end : std_logic;
        llr_mem_rd : std_logic;
        llr_mem_addr : row_addr_t;
        result_addr : row_addr_t;
        result_wr : std_logic;
        store_cn_wr : std_logic;
        store_cn_addr : col_addr_t;
        load_cn_rd : std_logic;
        load_cn_addr : col_addr_t;
        store_vn_wr : std_logic;
        store_vn_addr : row_addr_t;
        load_vn_rd : std_logic;
        load_vn_addr : row_addr_t;
        store_signs_wr : std_logic;
        store_signs_addr : signs_addr_t;
        load_signs_rd : std_logic;
        load_signs_addr : signs_addr_t;
        min_offset : min_id_t;
        roll : roll_t;
    end record;
function pack(int_in : inst_t) return std_logic_vector;
function unpack(int_in : std_logic_vector) return inst_t;
type inst_array_t is array(integer range <>) of vec_inst_t;
constant INSTRUCTIONS : inst_array_t(0 to 180-1) := (pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '0',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '0',load_signs_addr => "0000000", min_offset => "000", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '0',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '0',load_signs_addr => "0000000", min_offset => "000", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0000000", min_offset => "000", roll => "00000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0000001", min_offset => "000", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00101", store_signs_wr => '1',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0000010", min_offset => "000", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "0000001", load_signs_rd => '1',load_signs_addr => "0000011", min_offset => "001", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01011", store_signs_wr => '1',store_signs_addr => "0000010", load_signs_rd => '1',load_signs_addr => "0000100", min_offset => "010", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01100", store_signs_wr => '1',store_signs_addr => "0000011", load_signs_rd => '1',load_signs_addr => "0000101", min_offset => "011", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01101", store_signs_wr => '1',store_signs_addr => "0000100", load_signs_rd => '1',load_signs_addr => "0000110", min_offset => "100", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "0000101", load_signs_rd => '1',load_signs_addr => "0000111", min_offset => "101", roll => "00001")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00001", store_signs_wr => '1',store_signs_addr => "0000110", load_signs_rd => '1',load_signs_addr => "0001000", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '1',store_signs_addr => "0000111", load_signs_rd => '1',load_signs_addr => "0001001", min_offset => "000", roll => "10110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00110", store_signs_wr => '1',store_signs_addr => "0001000", load_signs_rd => '1',load_signs_addr => "0001010", min_offset => "001", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00111", store_signs_wr => '1',store_signs_addr => "0001001", load_signs_rd => '1',load_signs_addr => "0001011", min_offset => "010", roll => "10001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "0001010", load_signs_rd => '1',load_signs_addr => "0001100", min_offset => "011", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01101", store_signs_wr => '1',store_signs_addr => "0001011", load_signs_rd => '1',load_signs_addr => "0001101", min_offset => "100", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01110", store_signs_wr => '1',store_signs_addr => "0001100", load_signs_rd => '1',load_signs_addr => "0001110", min_offset => "101", roll => "01100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "0001101", load_signs_rd => '1',load_signs_addr => "0001111", min_offset => "110", roll => "00000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "0001", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00010", store_signs_wr => '1',store_signs_addr => "0001110", load_signs_rd => '1',load_signs_addr => "0010000", min_offset => "111", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '1',store_signs_addr => "0001111", load_signs_rd => '1',load_signs_addr => "0010001", min_offset => "000", roll => "00110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "0010000", load_signs_rd => '1',load_signs_addr => "0010010", min_offset => "001", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01010", store_signs_wr => '1',store_signs_addr => "0010001", load_signs_rd => '1',load_signs_addr => "0010011", min_offset => "010", roll => "01010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01110", store_signs_wr => '1',store_signs_addr => "0010010", load_signs_rd => '1',load_signs_addr => "0010100", min_offset => "011", roll => "11000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01111", store_signs_wr => '1',store_signs_addr => "0010011", load_signs_rd => '1',load_signs_addr => "0010101", min_offset => "100", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "0010100", load_signs_rd => '1',load_signs_addr => "0010110", min_offset => "101", roll => "00000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "0010", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00011", store_signs_wr => '1',store_signs_addr => "0010101", load_signs_rd => '1',load_signs_addr => "0010111", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '1',store_signs_addr => "0010110", load_signs_rd => '1',load_signs_addr => "0011000", min_offset => "000", roll => "00010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "0010111", load_signs_rd => '1',load_signs_addr => "0011001", min_offset => "001", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01001", store_signs_wr => '1',store_signs_addr => "0011000", load_signs_rd => '1',load_signs_addr => "0011010", min_offset => "010", roll => "10100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01111", store_signs_wr => '1',store_signs_addr => "0011001", load_signs_rd => '1',load_signs_addr => "0011011", min_offset => "011", roll => "11001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10000", store_signs_wr => '1',store_signs_addr => "0011010", load_signs_rd => '1',load_signs_addr => "0011100", min_offset => "100", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "0011011", load_signs_rd => '1',load_signs_addr => "0011101", min_offset => "101", roll => "00000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "0011", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '1',store_signs_addr => "0011100", load_signs_rd => '1',load_signs_addr => "0011110", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "0011101", load_signs_rd => '1',load_signs_addr => "0011111", min_offset => "000", roll => "10111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01010", store_signs_wr => '1',store_signs_addr => "0011110", load_signs_rd => '1',load_signs_addr => "0100000", min_offset => "001", roll => "00011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01011", store_signs_wr => '1',store_signs_addr => "0011111", load_signs_rd => '1',load_signs_addr => "0100001", min_offset => "010", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10000", store_signs_wr => '1',store_signs_addr => "0100000", load_signs_rd => '1',load_signs_addr => "0100010", min_offset => "011", roll => "01001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10001", store_signs_wr => '1',store_signs_addr => "0100001", load_signs_rd => '1',load_signs_addr => "0100011", min_offset => "100", roll => "01011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "0100010", load_signs_rd => '1',load_signs_addr => "0100100", min_offset => "101", roll => "00000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "0100", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00010", store_signs_wr => '1',store_signs_addr => "0100011", load_signs_rd => '1',load_signs_addr => "0100101", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00011", store_signs_wr => '1',store_signs_addr => "0100100", load_signs_rd => '1',load_signs_addr => "0100110", min_offset => "000", roll => "11000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '1',store_signs_addr => "0100101", load_signs_rd => '1',load_signs_addr => "0100111", min_offset => "001", roll => "10111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00110", store_signs_wr => '1',store_signs_addr => "0100110", load_signs_rd => '1',load_signs_addr => "0101000", min_offset => "010", roll => "00001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "0100111", load_signs_rd => '1',load_signs_addr => "0101001", min_offset => "011", roll => "10001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10001", store_signs_wr => '1',store_signs_addr => "0101000", load_signs_rd => '1',load_signs_addr => "0101010", min_offset => "100", roll => "00011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10010", store_signs_wr => '1',store_signs_addr => "0101001", load_signs_rd => '1',load_signs_addr => "0101011", min_offset => "101", roll => "01010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "0101010", load_signs_rd => '1',load_signs_addr => "0101100", min_offset => "110", roll => "00000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "0101", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '1',store_signs_addr => "0101011", load_signs_rd => '1',load_signs_addr => "0101101", min_offset => "111", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "0101100", load_signs_rd => '1',load_signs_addr => "0101110", min_offset => "000", roll => "11001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01001", store_signs_wr => '1',store_signs_addr => "0101101", load_signs_rd => '1',load_signs_addr => "0101111", min_offset => "001", roll => "01000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01100", store_signs_wr => '1',store_signs_addr => "0101110", load_signs_rd => '1',load_signs_addr => "0110000", min_offset => "010", roll => "00111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10010", store_signs_wr => '1',store_signs_addr => "0101111", load_signs_rd => '1',load_signs_addr => "0110001", min_offset => "011", roll => "10010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10011", store_signs_wr => '1',store_signs_addr => "0110000", load_signs_rd => '1',load_signs_addr => "0110010", min_offset => "100", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "0110001", load_signs_rd => '1',load_signs_addr => "0110011", min_offset => "101", roll => "00000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "0110", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00001", store_signs_wr => '1',store_signs_addr => "0110010", load_signs_rd => '1',load_signs_addr => "0110100", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '1',store_signs_addr => "0110011", load_signs_rd => '1',load_signs_addr => "0110101", min_offset => "000", roll => "01101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00110", store_signs_wr => '1',store_signs_addr => "0110100", load_signs_rd => '1',load_signs_addr => "0110110", min_offset => "001", roll => "11000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "0110101", load_signs_rd => '1',load_signs_addr => "0110111", min_offset => "010", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10011", store_signs_wr => '1',store_signs_addr => "0110110", load_signs_rd => '1',load_signs_addr => "0111000", min_offset => "011", roll => "01000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10100", store_signs_wr => '1',store_signs_addr => "0110111", load_signs_rd => '1',load_signs_addr => "0111001", min_offset => "100", roll => "00110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "0111000", load_signs_rd => '1',load_signs_addr => "0111010", min_offset => "101", roll => "00000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "0111", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00001", store_signs_wr => '1',store_signs_addr => "0111001", load_signs_rd => '1',load_signs_addr => "0111011", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00011", store_signs_wr => '1',store_signs_addr => "0111010", load_signs_rd => '1',load_signs_addr => "0111100", min_offset => "000", roll => "00111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '1',store_signs_addr => "0111011", load_signs_rd => '1',load_signs_addr => "0111101", min_offset => "001", roll => "10100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00101", store_signs_wr => '1',store_signs_addr => "0111100", load_signs_rd => '1',load_signs_addr => "0111110", min_offset => "010", roll => "10000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "0111101", load_signs_rd => '1',load_signs_addr => "0111111", min_offset => "011", roll => "10110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10100", store_signs_wr => '1',store_signs_addr => "0111110", load_signs_rd => '1',load_signs_addr => "1000000", min_offset => "100", roll => "01010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10101", store_signs_wr => '1',store_signs_addr => "0111111", load_signs_rd => '1',load_signs_addr => "1000001", min_offset => "101", roll => "10111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "1000000", load_signs_rd => '1',load_signs_addr => "1000010", min_offset => "110", roll => "00000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "1000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '1',store_signs_addr => "1000001", load_signs_rd => '1',load_signs_addr => "1000011", min_offset => "111", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "1000010", load_signs_rd => '1',load_signs_addr => "1000100", min_offset => "000", roll => "01011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01010", store_signs_wr => '1',store_signs_addr => "1000011", load_signs_rd => '1',load_signs_addr => "1000101", min_offset => "001", roll => "10011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01011", store_signs_wr => '1',store_signs_addr => "1000100", load_signs_rd => '1',load_signs_addr => "1000110", min_offset => "010", roll => "01101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10101", store_signs_wr => '1',store_signs_addr => "1000101", load_signs_rd => '1',load_signs_addr => "1000111", min_offset => "011", roll => "00011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10110", store_signs_wr => '1',store_signs_addr => "1000110", load_signs_rd => '1',load_signs_addr => "1001000", min_offset => "100", roll => "10001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "1000111", load_signs_rd => '1',load_signs_addr => "1001001", min_offset => "101", roll => "00000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "1001", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00010", store_signs_wr => '1',store_signs_addr => "1001000", load_signs_rd => '1',load_signs_addr => "1001010", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '1',store_signs_addr => "1001001", load_signs_rd => '1',load_signs_addr => "1001011", min_offset => "000", roll => "11001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00101", store_signs_wr => '1',store_signs_addr => "1001010", load_signs_rd => '1',load_signs_addr => "1001100", min_offset => "001", roll => "01000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00111", store_signs_wr => '1',store_signs_addr => "1001011", load_signs_rd => '1',load_signs_addr => "1001101", min_offset => "010", roll => "10111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "1001100", load_signs_rd => '1',load_signs_addr => "1001110", min_offset => "011", roll => "10010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10110", store_signs_wr => '1',store_signs_addr => "1001101", load_signs_rd => '1',load_signs_addr => "1001111", min_offset => "100", roll => "01110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10111", store_signs_wr => '1',store_signs_addr => "1001110", load_signs_rd => '1',load_signs_addr => "1010000", min_offset => "101", roll => "01001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "1001111", load_signs_rd => '1',load_signs_addr => "1010001", min_offset => "110", roll => "00000")),
pack((row_end => '1', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "1010", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00100", store_signs_wr => '1',store_signs_addr => "1010000", load_signs_rd => '1',load_signs_addr => "1010010", min_offset => "111", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "00111", store_signs_wr => '1',store_signs_addr => "1010001", load_signs_rd => '1',load_signs_addr => "1010011", min_offset => "000", roll => "00011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01000", store_signs_wr => '1',store_signs_addr => "1010010", load_signs_rd => '1',load_signs_addr => "1010100", min_offset => "001", roll => "10000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01001", store_signs_wr => '1',store_signs_addr => "1010011", load_signs_rd => '1',load_signs_addr => "1010101", min_offset => "010", roll => "00010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "01100", store_signs_wr => '1',store_signs_addr => "1010100", load_signs_rd => '1',load_signs_addr => "1010110", min_offset => "011", roll => "11001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '1',load_vn_addr => "10111", store_signs_wr => '1',store_signs_addr => "1010101", load_signs_rd => '1',load_signs_addr => "1010111", min_offset => "100", roll => "00101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "1010110", load_signs_rd => '1',load_signs_addr => "0000000", min_offset => "101", roll => "00001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '1',store_cn_addr => "1011", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '1',store_signs_addr => "1010111", load_signs_rd => '1',load_signs_addr => "0000111", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0001111", min_offset => "000", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0010110", min_offset => "000", roll => "10110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0011101", min_offset => "000", roll => "00110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0100100", min_offset => "000", roll => "00010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0101100", min_offset => "000", roll => "10111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0110011", min_offset => "000", roll => "11000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0111010", min_offset => "000", roll => "11001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1000010", min_offset => "000", roll => "01101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1001001", min_offset => "000", roll => "00111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "00001", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1010001", min_offset => "000", roll => "01011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0001000", min_offset => "000", roll => "11001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '1',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0110100", min_offset => "000", roll => "00011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "00010", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0111011", min_offset => "001", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "00001", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0010000", min_offset => "001", roll => "11000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '1',store_vn_addr => "00001", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0100101", min_offset => "001", roll => "10100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "00011", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1001010", min_offset => "001", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "00010", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0010111", min_offset => "001", roll => "10111")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '1',store_vn_addr => "00010", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0100110", min_offset => "001", roll => "01000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "00100", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0111100", min_offset => "001", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "00011", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0000001", min_offset => "010", roll => "00001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '1',store_vn_addr => "00011", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0001001", min_offset => "010", roll => "10000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0010001", min_offset => "001", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0011000", min_offset => "010", roll => "10001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0011110", min_offset => "010", roll => "01010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0100111", min_offset => "010", roll => "10100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0101101", min_offset => "001", roll => "00011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0110101", min_offset => "011", roll => "10001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0111101", min_offset => "001", roll => "01000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1000011", min_offset => "010", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1001011", min_offset => "011", roll => "10110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "00101", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1010010", min_offset => "001", roll => "10011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "00100", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0000010", min_offset => "010", roll => "10111")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '1',store_vn_addr => "00100", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0111110", min_offset => "001", roll => "10000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "00110", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1001100", min_offset => "010", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "00101", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0001010", min_offset => "100", roll => "01010")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '1',store_vn_addr => "00101", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0101000", min_offset => "011", roll => "10010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "00111", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0110110", min_offset => "011", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "00110", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0001011", min_offset => "100", roll => "00011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '1',store_vn_addr => "00110", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1001101", min_offset => "011", roll => "01000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "01000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1010011", min_offset => "100", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "00111", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0000011", min_offset => "100", roll => "01110")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '1',store_vn_addr => "00111", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0001100", min_offset => "010", roll => "00010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0010010", min_offset => "011", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0011001", min_offset => "101", roll => "01100")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0011111", min_offset => "011", roll => "11000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0101001", min_offset => "011", roll => "11001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0101110", min_offset => "010", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0110111", min_offset => "101", roll => "01010")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0111111", min_offset => "010", roll => "00111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1000100", min_offset => "100", roll => "00110")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1001110", min_offset => "101", roll => "10111")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "01001", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1010100", min_offset => "010", roll => "01101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "01000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0011010", min_offset => "101", roll => "01001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '1',store_vn_addr => "01000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0101111", min_offset => "011", roll => "11001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "01010", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1010101", min_offset => "100", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "01001", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0010011", min_offset => "011", roll => "10010")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '1',store_vn_addr => "01001", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0100000", min_offset => "100", roll => "00101")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "01011", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1000101", min_offset => "100", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "01010", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0000100", min_offset => "011", roll => "01001")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '1',store_vn_addr => "01010", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0100001", min_offset => "011", roll => "00011")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "01100", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1000110", min_offset => "100", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "01011", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0000101", min_offset => "100", roll => "01011")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '1',store_vn_addr => "01011", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0110000", min_offset => "100", roll => "10001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '1',llr_mem_addr => "01101", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1010110", min_offset => "101", roll => "00001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "01100", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0000110", min_offset => "100", roll => "00000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "01110", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '1',store_vn_addr => "01100", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0001101", min_offset => "101", roll => "00001")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "01101", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0001110", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "01111", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '1',store_vn_addr => "01101", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0010100", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "01110", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0010101", min_offset => "111", roll => "00000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "10000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '1',store_vn_addr => "01110", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0011011", min_offset => "101", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "01111", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0011", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0011100", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "10001", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '1',store_vn_addr => "01111", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0100010", min_offset => "101", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "10000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0100", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0100011", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "10010", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '1',store_vn_addr => "10000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0101010", min_offset => "101", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "10001", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0101", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0101011", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "10011", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '1',store_vn_addr => "10001", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0110001", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "10010", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0110", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0110010", min_offset => "111", roll => "00000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "10100", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '1',store_vn_addr => "10010", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0111000", min_offset => "101", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "10011", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "0111", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "0111001", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "10101", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '1',store_vn_addr => "10011", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1000000", min_offset => "101", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "10100", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1000001", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "10110", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '1',store_vn_addr => "10100", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1000111", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "10101", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1001", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1001000", min_offset => "111", roll => "00000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '1',llr_mem_addr => "10111", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '1',store_vn_addr => "10101", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1001111", min_offset => "101", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "10110", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1010", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1010000", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '1', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '1',load_cn_addr => "1011", store_vn_wr => '1',store_vn_addr => "10110", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '1',load_signs_addr => "1010111", min_offset => "110", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '1',result_addr => "10111", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '0',load_cn_addr => "0000", store_vn_wr => '0',store_vn_addr => "00000", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '0',load_signs_addr => "0000000", min_offset => "111", roll => "00000")),
pack((row_end => '0', col_end => '0', llr_mem_rd => '0',llr_mem_addr => "00000", result_wr => '0',result_addr => "00000", store_cn_wr => '0',store_cn_addr => "0000", load_cn_rd => '0',load_cn_addr => "0000", store_vn_wr => '1',store_vn_addr => "10111", load_vn_rd => '0',load_vn_addr => "00000", store_signs_wr => '0',store_signs_addr => "0000000", load_signs_rd => '0',load_signs_addr => "0000000", min_offset => "110", roll => "00000")));
end package;
package body common is
function pack(int_in : inst_t) return std_logic_vector is
variable rv : vec_inst_t;
begin
rv(1-1) := int_in.row_end;
rv(2-1) := int_in.col_end;
rv(3-1) := int_in.llr_mem_rd;
rv(8-1 downto 3) := std_logic_vector(int_in.llr_mem_addr);
rv(13-1 downto 8) := std_logic_vector(int_in.result_addr);
rv(14-1) := int_in.result_wr;
rv(15-1) := int_in.store_cn_wr;
rv(19-1 downto 15) := std_logic_vector(int_in.store_cn_addr);
rv(20-1) := int_in.load_cn_rd;
rv(24-1 downto 20) := std_logic_vector(int_in.load_cn_addr);
rv(25-1) := int_in.store_vn_wr;
rv(30-1 downto 25) := std_logic_vector(int_in.store_vn_addr);
rv(31-1) := int_in.load_vn_rd;
rv(36-1 downto 31) := std_logic_vector(int_in.load_vn_addr);
rv(37-1) := int_in.store_signs_wr;
rv(44-1 downto 37) := std_logic_vector(int_in.store_signs_addr);
rv(45-1) := int_in.load_signs_rd;
rv(52-1 downto 45) := std_logic_vector(int_in.load_signs_addr);
rv(55-1 downto 52) := std_logic_vector(int_in.min_offset);
rv(60-1 downto 55) := std_logic_vector(int_in.roll);
return rv;
end function;
function unpack(int_in : std_logic_vector) return inst_t is
variable rv : inst_t;
begin
rv.row_end:= (int_in(1-1));
rv.col_end:= (int_in(2-1));
rv.llr_mem_rd:= (int_in(3-1));
rv.llr_mem_addr:= unsigned(int_in(8-1 downto 3));
rv.result_addr:= unsigned(int_in(13-1 downto 8));
rv.result_wr:= (int_in(14-1));
rv.store_cn_wr:= (int_in(15-1));
rv.store_cn_addr:= unsigned(int_in(19-1 downto 15));
rv.load_cn_rd:= (int_in(20-1));
rv.load_cn_addr:= unsigned(int_in(24-1 downto 20));
rv.store_vn_wr:= (int_in(25-1));
rv.store_vn_addr:= unsigned(int_in(30-1 downto 25));
rv.load_vn_rd:= (int_in(31-1));
rv.load_vn_addr:= unsigned(int_in(36-1 downto 31));
rv.store_signs_wr:= (int_in(37-1));
rv.store_signs_addr:= unsigned(int_in(44-1 downto 37));
rv.load_signs_rd:= (int_in(45-1));
rv.load_signs_addr:= unsigned(int_in(52-1 downto 45));
rv.min_offset:= unsigned(int_in(55-1 downto 52));
rv.roll:= unsigned(int_in(60-1 downto 55));
return rv;
end function;
end package body;
